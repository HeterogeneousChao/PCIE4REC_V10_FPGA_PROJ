// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:19 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bsof+xwDQSfnlB7OyFpIn7y79oUC0VJFJZ8FWdG2l9Gkgk1vb4F3PQsPClE7TluV
2vGGa4VePnTiCC5fvAAqQqm9EPqbO6v3oEpOKJ3O3nxwX85lt6OVT2x7xfRTWFim
n1TWG+pvaJRZYW4/Lx6YDQVvi5Q3Y8osRBs2tiDQLZg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
9bXNwaelCjC01kthYrLDnl/WMT7LDUgby3cojindKrNAYJSCsdMrW4CLlBn4NJXK
tmLP2hdWwI+ZME+1SvFwCw8VADGg/1JgOERuBPumFzLI5xldbF45I1Ij1vd/n3KY
s6AP+qyLk9CJz3VoR0TE7ZRgmoE+KFVxmBLFrDFyH6zQ8it9a3OaB5HvAYQCVkbl
HCtqylKmxsik3Wr7G9gtGcZZ2+gg7teNQoMJI5FHGPOaI/iPdwpKzcYU6tqWWTGX
xUkVExZltwGQ3a9AON/ocwOWLxEXrfKnalahWWciKhOT8ZgpUMIYtpG8Mw6rVJXS
9orsHYt+tEwLOuCIJ0jLsxVxCifJ4QFobde7CoS8TWMJiWoQh5posoGzhQ1dfyMO
sJxG0dZMLqjh/UPSHwssWTReP/xZiWxkTYVQHxrJOmb9yB9SmsaqG3DGXTYFZEAc
BDNSvOKcI01I4wngdLTofkJzRqW6qBMBN8D2G+A+FyWQPRi/XKuZSLKEMy0jkPlE
pYLM5HDMHa6SnCrBW7hUOOxsRAgtYOrSgoytC7gWCcdYboegdn/0MC75+FswSAyN
fmGJxuXHBFBcnu4ij/xmxryRFEFY5Y6bPTlHxXNFUIWK25qTWWQsxFRQAk2kC362
i30sMPxTleGVKUS57I2JU4gtKhVSywYTAE8rGuaKIIQKkofnmmrrnpPCsGFjsDgv
DYQQC7sA2++gKtW0Bd5zw3EWiobwYk9+XC6h/ZrzpIrD+Mq2v5OgWaRS+kWaeTet
3h2hpeba6hMvjQ4nx8r7uTzGSV9OyeWKvSerUR4uIyQEq/PAaA7lJso4N8idipPw
WkxfsL1oH16IlgQj1tjsBKRKoHtmnabLsaqC5cd9jeJLZpM+pLTfukt9xgS+k8cP
O37tIy5yROLfjv+cZSAA4RW1DRBeUH/FfdsKL3xE8XFhpi0GaKmCRahSHV4fyR3u
QB3BZF4+0BITeaZ7BwrjqhpA+oerME8HHgwZ1RXv4VV/zEAV9idU7DzMpKxXlIuE
aC//woKCTMquT4TjbquPfMVj4KG0B1GStWVml0RDQcX57ZL6OUgKeaMumvyLhyEf
gh3TUDDc8oVL1SiFk5/BOM/WswUUycrXhQ1/y/hkghzcF1Xt4v5Qu/h0sOA+pb5f
2qZzkm+YWRXIjSZ3cI7mQSiPMKE7Jfv86aJ9PRa0FwiM9+1UN5ImYhzigHZJDNmo
/ORj4t1jT1yCHjHDP7UuSh6UwcUlOSpZJg+faJlpPlISZBN9HLr3uOiYCYPka/Ke
t78g1omUgmwS2mNSoTYhQyL33/Ofy3XPniCQPoHORzNS6rkXdW0+DrMjWGga+3GM
PDqgWirg8fDN6MvrlXZ/nQWvM0ysICfl0PT23p89ytWzLPl13YmH/AeZnGI+Y7Ac
2kcIJdTTBdDRLKGu21bF3ADRh1oDDbERdA8aGTEK3ukmmUwdwQKHJ3ZGQcjY2e8R
Iq6J1veDRB3iHGYrGahfk8q65WBKTUNzNj/lPzNgFpLaPgYIo4GIjBBPF2YIdUzd
x3VEa766WNoyLzlCpMhJEqxwf8Ogv+jLBSwXuAP6YhCQWeqTh0C5Iy5MlkBDx/cU
22ANncj9pXRWdQrhv2C49WdIF6ZZnsIYN+fkerLhJn675dw/eoVlwQLb9vaiw99v
KVquXoCQKQV9aVRmBXzKPsI2/i9lLXAZf9sqqA1oj4/btO24WWzZdw0BL91KoEtN
l7FFEaGwAV79WrcPs3zKq7IUr8A69ImHROlcvgeZIqycIIh0f0TZFpQXOrMUAhRi
HVa/mRiwsLCpDuGs6sBDvFDWpgdTYuwx0lIUkc3TWPI2ILcrLKPb6P1cPZbugo5y
KkR28Qjj5bDOJ7GTLq5O99q8uV4J6DY1dE1zHN9fNySLPpbKKP//kF+mZXodDIS7
UGYtOn7enHxIvVVj9AYOxRlg0nglaxFSJKmS5QaEbZG2lOD79UPwerylYBcxcz0e
+LQB7YjeARD8AYwiasKYjshZMAPxyvBDEMKWKybl5TEgo9CxuJsQs656kcDMWr6z
RTfHHZy9vkg2RB+r1oSdpuTH9z+gbgmgPUWfNkxMNzb9Rew+HOsjKyGlraUXCx8Z
i7k/xNM/qf1zuXZJYqf0VCi6yi3LwloeGgToTiUiGcD4cndby6+pGOg7RghqFYkj
zSMbhKCpArwFSvmpT3gbgH59nVzViDBfGJLmI6Enw9cD32X9u4m6q0D63o/qRQZh
uch9RCV4vLnyyqPyXTZGF3LlpnuT/IkL6lVBmBs7j3N14BBiUh8xu3xLv/IbtdaC
B7spiZC9CkSZBQa6GO/F2JvPFp/FypGtzceXOElAqSumRasrW1KqEBRye3dUhgIV
UC/SZu45DLf5t33rR8cVL03Uw2xoNKtj+uye0IVQtz7lxtaqoK0R+slncFk0zp/x
OJrxwsUWxTnJX45fiyyh06VmTy8yNcuuS4k4n/0zxrt2D7Q2IYXNOpBlJ/VOYIPX
J6xQXHfQ938wEL4cbndh+Axbf0USXe16rXys+QFVjTsnO1FZ/t38fRPH53152bGZ
e4weRboYsY7Svh/4KpEkPAjH4NZ03fdXfWntRja4adP5/6KkUyThkj93+HfohfmP
eTKrJuwnU4/AOWJ3O8nYFyusHv0JP48yGseuqCA2jS8mgLkG+cD7ePVKUcOif7nJ
s0OZgIdOQCXRQKNQ/r3PULgxXtCZwDpGwLSxKoPv22LmN8c/fWAPOSGcFZemYmtE
vGdLhQR/Qhw9PzrtGu9UdCAIVVrBEnPzuDXbgiTbGpUqH0FdzsmRhXylQbXUJUC4
yAswTDcxZAh88Y8y+X3YYvC8w2dEyN6Z/OW7qbQKajhYRgEytI8k+bxvlzywzPoy
iBPCIrOA9ejs0dMzf7CpzlMmSUIXf6bAjDfpYqF2ieO7bi4zDNIxNmZL08Zwe5Jv
sM/mdV/Tj+O+gFheZ57QoQ==
`pragma protect end_protected
