// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LkiCWIuBjNo2YTpm/rU+pAqNoEab+V6PPLvvXdvNa5yP2fHiYbYleFbbZB1EVdXJ
rJuCBpq0dtBh26AFCB3zfZEAj4+ZdHsUSeyOUKz8svEfHeZxAS5wuK6CRG9zZhJe
202d5Jlwi67jBKp6tAHJX+6P9WasIJUvckEVgGWqYQk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
VMMCStX8CdoWxBFhuXKHs4zvKaknovwphYQ5D7kRoOBtzb8m9ZWXLqfgr5lGMu76
bUW9r2D5tBrhUTmUnr1v/FF0TQHo0ufZwLyjNKVi+Y8UnjskLYL3W1TwLjxt19dn
SuHEOi+kq0itEh53YOqTfN4bq0zHTG3ca/KyTxUY1/zpLmHWUJmrAFmwM6LG4EXZ
gBWwuuHL8DQaEt6z3EqROhYbc4Q9NFm0jYcEa3EO39VUu8i5iMk+wWZdG6JqMv/H
9tAD9Mvci5fkAMEWiPmU/hFOY+ct1f/a1Lzsl99pGBt4T3JIqYf7NiMdnyMkO0DS
ObEUpZmumxyexikK2teeGkpex/APCsDHtzx/zply8ZZNfNEm3TxmmJS13VDJ1pVF
L8Fq6dua9DULgH77Yt1Sbh07rlfyNkmMjgNNFX87nvq99DXMA4YdET/SpS65gXqZ
8A/LJksBLZLot+KIp86MpQl6XX59UPecyPnmmMfi/B2aaHCU2fx6jWCRqRzcefub
B8O7cYdg07uEs5ppcE9zMocrwy0qUVhay3jwCP929AWO0vsxTzYHsxljpdqZ4AoM
Ac0ESK60xXm0EuGnjQEeGvx0lZ77rfwIJv5rQxXhcwAAEEn8lmkEvd0nKvSN3ujf
bWVqu0PPWbwNC06FKvg6VX2ZIncKoSOKySE2pPdRJ1jGYMMSwWlQarhKJIaVTaMc
L1TCYYJ/1FOBtX/wsxduTmjjaTgjuOxNpPsjHy1vgHF9ha/IQD/NfHhvExDjFKpS
yKBIYOcv/l7yWz5hLbip4IAS5RhJa6zplCurHhVP9mz6qIYRK6dw2eSL6LvRroDd
3mc91We+jiMFbARz2xHMjFKeO5l4ris9Ihl9bdqgpY32+RS0Y38WpapfhWkkb91s
aUZJwx5U6awMz9+b6FUqDET2rCG5Cez/mNGZ60Q1yJOXI+s3l3LOKh3jwTObwqPy
WW0wXysq2D4r5KGQYMDA15E5EFoz8yJjikGZmYYa7bRWDoIFFDAShm+PEgZm4cc6
GiqN7g908/jJyxgbzDSpAUaXtpdOP8B4/TcoAWNuiOIOAZj/rMu5otpnJ4sXRjRC
SNXIxkZVRSer+Af54HOytZqs4n6MPPlA82Ch71IjKbMs/Fk0TQWJj02z8y7TuNNC
rg4i7q4EtoOcQyoUxqbFDU4Ong1BvnmxtcBajfR2yvueqMXpgRpg58VyXJggMT3o
odaKSlSvBf7WdOp4kGj4iN6+Gssn6Dn1qCfl8EBw+grWSbHFAUgGnUO/JwmyRjL+
/G5xjlGY5hlV6iP/HacnF1Ou3I9qmwKhibPyUKjrgyYdyCdeQ6PiAVeCW3BI9wLS
vMbXOjiTNqtVduPBhwsTFEWZL5h8gJNJ3VIrKaJFPiuC6Ue2V2jT0CIDY79RE3+I
GGD6gbiJ5uNd1QowPJVN7uGpOAQCa35lnQ1IXDup3cR2xNCaCd9lbHMu/1Gxirb2
9O/ULu/LVfB0i4nbxeR5H5a64ANtdokO8GJlp+ybzZnB0W2r6lEdwVLdidlUm/mD
CJsf3v+i/9D9MrajISHkXX95Clh+8aXs1wFIkg/VxogB07tqkSayFiYQLnswPG5b
CV4xZIroMI8y7h0bZGlfb/UbiHTbQ4IEqu9gSjuwfU+qz4Hv2fqr0XvaJCxuw0Wx
8gxWnmpGBvtEncaBH3Zjxg+Jqrh+HAcy1tRhi4h8bD1+NabslS8F/UNxErTeMOOO
yIAeu0/Ewm1xzNE/mLTDBhdj+4Lig3+MLkT5Y7y8ym6hp3xSkDajoLmTx9GsH6kc
IDEEUKxSe3L8iwaxvoMx7zqDI7ozwioZUKu7XDKXgnm2puqUzzeV1dfQWZ6Jt4lc
YbAlb5KEgl/34wUtgVC7jHbC7fjzs6KfANPOu7Xjgx6DTwGmZDRpcGUFHWIZT3K7
jqmkEzM8uKrr81eK73R3lqbL/ZM1k+BX+fA0S7H4ZHe/2YK0gtvqdNIIBHfLrpm1
NiOS4AUpg4XbMPkrS7EeQt4cXw3xfXv4ufoXdficlUuGSEldNT6MhMo+tM3QodnM
E+Z9K7Og5nWx/1JXseNAq/sGy8z+fTOPcCfPaKGsvf9150P9EOQ5MViK37ixPb69
6S3SUtmTJ81K0jNGrFL+JvKpaPWUqZEBcKPBufoc36MwEk+4mGDPY7zN5S9Sxi1n
Zo32LlTWi8YKwif3Q4oj4XkywhrXc/+xCqYe8xotqlm5xnZ4EpK47jSLIsGczjGf
l88YhPLfjefEjR8LVko5Iiyutqyl1wZQKgFpMBEo7I67E3K/iIB0aozifi+7ETL6
a7AhauwOm47fuL3dn6xkDMmMKJmpduQ9sJbqDPITW7mfCMoAmQuI0I9XC01GyM9C
9h0whO+cBYs54lN76+MxVZegjcqxkAKCRSxpELTXjM4/KrxK4sMQh/oYpjS8s/DO
y8AZDo8TUIsaokGd/iCeOV2L+TpbiLMhCZqeIpq9WGu8T9T4nI2WEVfZVA2W59ST
gUVfhjOwGZNOzrW2VMP3bwYRSU7UXUuZCqKC7yHTTWb1Qoc/A7IBNCbeTNvP7rEh
IylBcVgAj5wrsWYGlvlk8OQ53lFi/2zj86VRkKa5kuRz2MSJxzYHVD8crtclJaS3
p0oh2xxa6A+fadHco0UtMsbS+YZ9nu6W2SubXKCfQGOB666YGdbo8/LO+BUtCyHw
boI+1Vt8BuyDidV9tJruMy+SjtduA5cHJA246Nr+z08Omj3zmUP6CxvvYmidDG69
Pcc0V/5QwOfc5c2PAR04Pox+e0ItZL38guJChCsiGWmjUZol986HQ1UNo7RrGBSY
pwMJO87LKK6UmsLKmeIbZk0SrVCoR2UsnNot6wkCoplwDLP1f8+yrbADb5vL+332
gLIgto8IP/bRPl1u0VRnj9GidUzp9cW8z1l0xk4xVmsfrKmSiqAGVD5HAJhnWpBz
fNqPWDPLmY8Gk7JrnUYQ34rlfsNFj77wK6lz2LS28Mi4RF6rc2Ev4tR6dQhJMozh
ymR76OGu0TQHu4+OtvyhDRZ3Yon+ql1e/RNp1rSFZmsoZtcEZ9ANKXKqJgsFrxj0
F/8s9i3UpEt0dQIhEngUxGkEBzTENBTvFd2Wgw5tbYvL5sgbmcD24t6/zV0Aa7KO
`pragma protect end_protected
