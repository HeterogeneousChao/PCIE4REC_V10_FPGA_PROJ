library verilog;
use verilog.vl_types.all;
entity DDC_1CHANNEL_SIM_vlg_tst is
    generic(
        clk_period      : integer := 10;
        clk_half_period : vl_notype;
        clk_period_1M   : vl_notype;
        clk_half_period_1M: vl_notype;
        data_num        : integer := 200000;
        initial_config_time: integer := 4000;
        time_sim        : vl_notype;
        clk_period_data_in_valid_low: vl_notype;
        INPUT_WIDTH     : integer := 16;
        OUTPUT_WIDTH    : integer := 24;
        CONFIG_WIDTH    : integer := 32;
        QMIXER_CONFIG_DATA_NUM: integer := 2;
        CIC1_CONFIG_DATA_NUM: integer := 3;
        CICC1_CONFIG_DATA_NUM: integer := 259;
        CIC2_CONFIG_DATA_NUM: integer := 3;
        CICC2_CONFIG_DATA_NUM: integer := 259;
        MHBF_CONFIG_DATA_NUM: integer := 176;
        DFIR_CONFIG_DATA_NUM: integer := 516;
        CIC_CICC1_CONFIG_DATA_NUM: vl_notype;
        CIC_CICC2_CONFIG_DATA_NUM: vl_notype;
        CONFIG_NUM      : vl_notype
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of clk_period : constant is 1;
    attribute mti_svvh_generic_type of clk_half_period : constant is 3;
    attribute mti_svvh_generic_type of clk_period_1M : constant is 3;
    attribute mti_svvh_generic_type of clk_half_period_1M : constant is 3;
    attribute mti_svvh_generic_type of data_num : constant is 1;
    attribute mti_svvh_generic_type of initial_config_time : constant is 1;
    attribute mti_svvh_generic_type of time_sim : constant is 3;
    attribute mti_svvh_generic_type of clk_period_data_in_valid_low : constant is 3;
    attribute mti_svvh_generic_type of INPUT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of OUTPUT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CONFIG_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of QMIXER_CONFIG_DATA_NUM : constant is 1;
    attribute mti_svvh_generic_type of CIC1_CONFIG_DATA_NUM : constant is 1;
    attribute mti_svvh_generic_type of CICC1_CONFIG_DATA_NUM : constant is 1;
    attribute mti_svvh_generic_type of CIC2_CONFIG_DATA_NUM : constant is 1;
    attribute mti_svvh_generic_type of CICC2_CONFIG_DATA_NUM : constant is 1;
    attribute mti_svvh_generic_type of MHBF_CONFIG_DATA_NUM : constant is 1;
    attribute mti_svvh_generic_type of DFIR_CONFIG_DATA_NUM : constant is 1;
    attribute mti_svvh_generic_type of CIC_CICC1_CONFIG_DATA_NUM : constant is 3;
    attribute mti_svvh_generic_type of CIC_CICC2_CONFIG_DATA_NUM : constant is 3;
    attribute mti_svvh_generic_type of CONFIG_NUM : constant is 3;
end DDC_1CHANNEL_SIM_vlg_tst;
