// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:18 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VTaEib+4N2WgvmJftivw8R6k6gnJsW7g1xT/wpAZ43tW+mfAzn0Fmx8hWOrTVpFK
JiURQS2/ITJ9VEi7d4D1tpGfiFpvWY1F45C+LihAHZFn+OmHMUifNZHKGaaFUZJS
FMKppsd3n+bhvHVOcLgHN0HjT58krSqHc5T9MpoJbC8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
H8EKsXjdDazf73TW1aNcE9pIKu5N9I3RsJl658xZ7QPY9sybjcEgN0hZP5uRVosC
M93mAaAIcXoUWptJByAseuXyXyJXHT+E8WTNk7PjF2/VWfc2Ufen/HLyomFnAckr
+HK3vpGFdHdWBHGsEOf1XTowwxVkW2smGiGPBc8qv4gHKzGeD4H+VWLuzlVad8oq
eLTTw9qA5HXEoZ6L48vRfl+6a1fr6KsFP5H5c23nIC4aeMDrUtdZH5NK1VRKcZDT
jh9OjjUcvXXMOQ4Yq0Q2i8vjpIHmDGPvNOs5XrcZfGeAIumjWgjNsE5Wyy3d+Jvd
bl9YWcb8c6Kfd1SUL5JFlq7FYHXf6sxYtH9IWDlMcTb3R16SLASb25IVCM5+QOLU
FUCTX7mLcQs1HeSy2PKM9RcOWwRZ6xLxX4EEQPVcsNibAhgF4T1svdtszet2MUpF
7DArAbKa+bL95XvOFmv6Hw3hviQ+7DpsQXnt3EWoXh1q3fx/XP57w8mytf1nconQ
4Pa1ApiJ8MdaTEj9OF1Vh7Srl0bxUmQgFKNGZ5XFgpyorzKzJs+bZDZpfoaGGe2O
M5o4OzXs5v4YnNjcNDr5Gyh+uZ2rZ4Fyzwa7UyppiCbaLeIzX0Dwosvx1tOg542R
1vIZJjpMWy3Q2C17WkuRqJUA5EgS4y3+Bo/zJXcx0T2MlNBmHWlVKFXlsVHk4p8s
Abk1fq2HvKOHvuoN5gcOmR6bpmMwSahYrPozvydWkgpHk9T68ktyLa+CRtBm6tBJ
EmDohVcv4lO78LomJ2NImWbRNgSIKWTB/JaBoTBSsnZifL2tGPN5t+yLOwpuW5fE
Swlwhv20CLEyj1P//ql0t9F4aaTy7wGlhV+FIzm9srffIrBnxdrg4jXgaZlmD5jP
NazJlmJhyXV5kMgj4sxdERwHv5vc+yY+7bAsFTdgABtlOhjeUNVW14IYLirhXIOt
adVvBpFpzYqdfzdHhMinTGBF3bfYhDHKL9EBpcby0LYIlwvX94zyqDHRpRlVssV9
js1Lfk8yzvpM8uFm1MyGBfhQdtJy0zGO2AyvNvcMJHhzneI9XVi/nVzplw6P7GOk
Fv+GFJRcGGqQKR6XnXElLW53guu32uS44V8SkUuErPSHFZMEkQiDI3YmLw97cn2W
kXdzVoa15TVhRLkQLRgNHb3xErB72Is+wJOe7GrRuH6irnQDEtp/jtLJ/08q2qdh
16rM7MruOJQpWMWU/VjzGIsrMLrXNZ4pT8FNpIRCGcV7A5car9uW939FQbgbkQxS
c5Gjw7S3Q1YrZf146RxlUzJiucR8+n6Qh7EBP2PK8+s/J2DvnD1Xgu4NuLqFH8eD
rZaeR/6ViAfAnWx0vwwcOOmK3oLmlccSpUZxVHOCI4yRTUymb2oGY0b8YED6vfcQ
/8Lu8MzeFNXn2FWy2C9uQP6IeyunWn1mFW0TCuq1LJ/mZyZtdKgtQ8/Egwj9nGdN
kuwxAIvmMoULthzrtVZXu4rO8Y4Aj7fT7xqmFQTnnkNpkKI9hvzBZySi1F82M53r
QWxCtRECgJnDumD3WPvZHf3Qa0qpGfbBBebMwG4ftUKiJ0Yu3VzZdnQTdFVgziYB
7RbH0zmFPK4mLAXHsjLX3pcNBH38ofPmN8+xKSCorYKJeWj3o4qZ5pMBjQPRsSwt
K4Pom3keFLjJBnQz2ES5ShnYAZG2iqWVm9h3srRNn2D5HnJ7N5RL0bV9yE5KGAYs
R20DzGWLdCCwCB0BCg0ZQ7AlMTQgzFb1kwvk0bETZpyBCl41rlm35HEcLpeAkvKZ
FCIKzYk+QDYYjsC+a3VZqozhJXq/L17CnCABUK8AB4BhDcDzLyEsubY/vqhycZ58
JiJT2DuMgmTrn3m8zQP1FlUrHJcifFD1KV157xfDdbMFNOBP5FxR5IIC52LsZgVT
ADAll7Z4fyjMvW+ntdHR/eReRkT7mHdCb7u0XTiwyH79vZ3LoCOdquWalgsqzz/o
z1RMaraD4364VldUM6gq9q9raODvFxrFhcOsjtNaCHfCaGqCbVCxUkhCyUmX7dsJ
FEkiZivnXRVYKVLNSYTJWp+cqI6V1UfXXpwbh479Hoq1Vh6btBgA/ZwcS4orC6Ww
3VwTYi7s8Larxw0c+fvLW9hddBd9PibQfjGqMk4/r03Ys2I9SdL+1EJXxkVqATum
3+lHmRDjr6HGkj38H7BPjQ4MBycYtLkfhXxP5IFmh2Qwkbl4iqU3jWDuXkjg3QHC
dNXecUxqkzrgoDjpDkPOcZzs9JeJnj9rw+TZO5RIe2fRK6V67FxINlU1yqOUQCk0
+2/f+zNXl/VH4HTWl3ImoC658rMR+NYSlMcyW5YcN++1nxmLNvf1UHrKZjc2K1rj
aoxhp0IQszLoj/l9v4HLweInbg6AXP8xam+T6f+OzG4BWaBbjpcDmCJT9Km/Hmfd
2TVM2Q+jGadKpRtOOsne+rQezl52Kh8NwW1gaxfCS+G0hLrp8LUV3EM1vrLhxEaZ
LpROa2f7crue98SneZo4t1a8Md3rSYL42KlRPTgn4+b+mGiVx3cZa5sWuUD21Ubj
CuiGiSzAKJIZ9EIhIE3NVgk9S5ma2/Q85amR4/jyrmP2vgV8VDi/E4ISH04s8k65
gYzBOlxEDBnD2rVKjkreIWLbCYyfl88jqeXNGr8CFQXopOg0X4ek/gP17Ray3XF3
zJwBySCtC0lXSG4T1L/+CXUPtJWw4UILasoO6uA/VD3O7C11wUjs44GSjC0xPPrx
hqYvXZi6ZB158sUbtZh8HfDsyIUttfUdnmqfwp4cQznDSy0Jt5dgeKw93EYWPXGX
YuIZiXeW2pfQuMU5ipIC6ZnomedvIGSdbMjSpKKde8Osat41ON4qzT5+oZcFJe1I
nqrWX3FXbNA3qpgGbgxr+HK0jUFl7QFYMx7WJkZF2HqLmUxyM5qJ3mJRPpJzhL3v
hZXv8vogEBUCD04erzT+ZvarRFoueEk0Y6bG5+DTGmtFK8s7XdAaWCLpLzClsKPR
i3+44muBQmhy5mCA1xGUnZbU7PzTM4DzajoyRyi1XoLaKmeWx5qmV6GuxhXdddyH
Vop4o6R3pjxwGdhnTu35fkSUv2m8SIhXujC0O05jTXZHRLA0sZSKN6Q4gAquJhtD
N6eVWbyMaxSQVaMpCmYzs/JAp/ZPIt5jCcQn/sengDTie6f56KpNkqmy/Tg7q81g
rRBPSqwurX/37CmaVL1i1BxU5xilKeEJWQYjghIeIUH00Q1mybTWe4xLsoCLw1hc
cZEwK94gNfYgx3meMqJqx6pMnodKjDqJHsotLQ7FMofRe6bOib5YuBzrVRJb/xul
HTriyer6hfKznRQYr74H9tsK7cwK+ekFvAxSCCbqOcjXxNDt459Ut1PC+tfOw5AV
c8HFym1xbpCahiHwrZ05KeouN16C6dGK3O6sgUPOpIbgAfjGdl5U5qEw8tC7bv1o
CicgArLdDFZiJSto8zgAsGIEzBLeMsltSlWcMHhd/GyrYJT2wfDqqMLkUyolcusO
s9dU1071/F46sYgTU5YLHRi3Vb1uO3jIdCEzsWvlzlWYismHiNFWL3FtzcFNTQm5
6u5Zlidop4VVJBs8S56p3tGWinYI9NfDdrVVHrTN1LOSRr0VQoVzZqDj+1yEE0gZ
plpnseBd301una0vRnnmN16dHdDi+Ny3tas3R6vO6SbZ4k1xpOTOXbQsNwXJPS34
2b5xosCo4aIrQTco5ukhlAbJByV/gy5yiJR7ZY9LF19q9x3eXCbF91nNecMKGD3C
Hg7zNEH2GzCBh1IzM/D4EWa83OBlbug6589l6Zzi3ZmIqFYMKPbemE3oXLYB6N8h
83ZVE8Z8kWL1juckZgxM3yg/QGCra6oj7kN8wVPvCVnc/7GS0jzyRhIrxsiTWkB+
STNSjHh9Aj+DODdMIv/iDcr3nxJg5CcAeQIOjHLBcT/TdgAdodRFtmgxw955E77W
XIXzP3lqBBgr6NKoEqb3uHN+KtEXwC/0OgSRDvpxd6A24EG093KIUhlJrFfW4DLe
mBI6lWtr5cXM1b7ZWEqOOrKPc7QSTNJX7VflgZJcJyqk29hMaZOPOrUlmeMM2M7P
JQSNv5UczmazFPNtwZD3CNr48f1xtv7dpR2Dnj0JQ6owMOIsRXgQQpOoiyTyhkp3
pnqTTYp6m6mUPG2M1WO7HcqNbk0Fn69h9eMBe6Id32BvVl/h352PNre3CkHT4ysY
aGXyqjOW5S3MnHXUo5hjtLsGKp9QaQL7Sp7jErnpFufNkEI7KLulimhG1V8JXsuI
C24CjJkgjell9iOlLdKTlRuHRnu27C2UVxwaH1lUzeIArShg9KPpGsjGH79hoBIf
Cv0o+/8TflfMiqPS2hHulg==
`pragma protect end_protected
