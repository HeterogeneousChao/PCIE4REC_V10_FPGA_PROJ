// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:26 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RBy5/YFow1XmyapT/ch2XJWQZvs7lXWb7XJWeJwCVZadapzRYWihqHV9zu+OrJA6
v9HnNbS00HNdMdFsw3Hs9yWExRT5X9Y+tkTDnrQY+I2z94ITJM/vzz9poueBL43y
q+3TBDGbTuvoXgcV9JtgZXdgR171irbnbZxS3AOe0SI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20992)
YKx8Fn5xhF6rGN/uI/odCAD0B7Bkxz/e8juUoJ1jwvGNT6yCQpZuU17omNyq6EcH
3bEuvyq2kJpOBbVpBKJ1WPzcOVvt/w1SeH6zQP+ZSfHD42eUCXm0LfpR0feSkjQK
1BHCJf4A5aDav3Fa1a/xK1rqgMqdGkIezhaMxy4KgSIE7hQnXUVi1gGODs0xphen
wh3KCvUMfc7Mm/jeJ0iML5lCjCmHkGGohwWBHQ8pOAeArAdr5O38t7K+NK3ZK73e
FgrXEOaW9S2GkY3gnWPJVwOoKELu0RZotsmUQJghDZe0XWvc5056vv5oBLGGxZBp
58uuVRYFT30aMC0sqCZr8F3TJlWlmosg6crvYPP483V5bjHoITIJjdPh8YMumuQe
31JNJznwGhHvfk8rr9yrhb0yabiNwhFGnmBQ+GUIj1XeAhDLOY4PT3JY6neVaW6W
WRQ3zF5CvAp1UZWA80fWH2YFkDNZTkhtprUe1lVEgEcy3uh8kwstqqRnIBrX+cE4
POB+RuFDOY0sX5x0i4QaWfqXfIQCpwSORYMVYfafS3xxGGMVEUwYCMuryrUKMc5J
PnfqVLOYdDBlQAb9DDUY0zx8fE+AUFEXYWJ3JDlcoWZTe/6TVO7c5yW98fqJ6JgT
TxIRT8kJfHsG0FC7wzmL1ePwz4FKCEGTf4be6Ps5m0BVRbvfB9oLl0o+ufTveAjs
CkqRBIPZms5gu+bFCeO1xynn2zBUgW7SUukBriOPpyeidJljbo1LqHELP0cRZxXX
HK5Cd2khwLDl0nke4Ekla70071h6oaBsltWG8RxymD+soSYqavHkrvO1Jtiqovg+
78KrD5uwSKBofIe5wNH7R0uZrFMTRw6VgqwWNr7Bqqav/0qLtSSwk3kqgvz7KC5C
jpVC+BN+UHFRDtEoSLWdxKH5Xkxh9a1E/uspFeiibQA3fl+4wB1oYlVdm4cpJOaz
pjal321/kniEqBSkyzVj3tJDXfy/ltbmeIGUKVY83hOCoxY2Nbpd+8TxUC1aCtmZ
29xin+A97Yt1Pe3gfi1xHMKcVFjzoP4HD0miO2HH2gcGsmV7j8ZGJipkTpiUNvRJ
N3UT2H7hM3Nz6poWvrxKk6rqcB9zJ3bUr8afoX2Q0/bQbjLeZVXUtSBRpFav8ZDd
Y3Oqz4h9unu07EH82hwYkdgacTjBC096hLZWM8HMGTtI3iZBl1JPqJKJu6lh7ar/
cJhY1fgBMsiVS1MvQoH+XXZ1iTx6hMAn/94Fr3h0EVCn1kacx5+x9A5wZbS/Glmt
h37vda1NKGijkY90IBCLIvbCb+8tjt4ip4pIrli0BXVHiwQZv/diVsDN/VyCKCaL
rf7n01umFhyhOqHd1d9AqZIZLL2tV88oLrV6N2B9u1t+zyLKYSaaZBTQoqIiAGAp
EPdZy7T0vg0kXUnj25MPsiG38ohRWiMAK2Q38sl9xiXGVBQIizR7atn4Pda08miH
BiPUF+GRAbz2Cl/FdzxuL6o+piSztCfWmTCQfVSHU7v2Kh/1+X3AIxeMm+gBI4H6
8VoB8Q4gqoTWuYCSXwUqeG23k3Fmx+BXD5hlhNsqCCEk0asLMdKbKrM08buNqQlv
3Bjq/PSR6+sJqG83u3SBZqicTOczDzHvWOjIScSh7Zm9xaGef9TKfn4piPoG8+QT
4JqGpwLZptvSu29pSglHhwJqLXTRkRigGVesXqILfjfkQS+Wv9pQKx2KLhUflORR
KwzEk4GCdEJbcoJMtJjEy4bZ88zYlcrDXU93TKCeb45OM2XCB2DNmAH5FOryh/XW
laYnidBYmGnraRuGXyQgJlAXsWWwK5Sn0+TcyNUk2ZCBt4HaiUrqPZjyIhtt++Bz
caUPAc22TRWCexKKcBWprSJo88d+Hl0iA8s9M0F3jFIvVOX0ZMtLmOoeQi+RGBiO
1ko8EwPqn17KJFWpxkk01Sj37xqkpiQa/i/hWGS0zAFG9jlcf4zmgy0eBHkNZzBm
ZKB7FXD+z5tUMwULJYqyUWboP8G37elUgnrfjbSFMNaSF+nIXpUnn3n9WPIbLLvb
3sz9HlAbYMVWrFtg0mnawF/n6eiH+0hsP9PNHgP49nNK4aohjahTJIbl9+CnFaz4
OqL78JcttQIX0z5i2Buva2ZWs7A7fz0J6BBuswyP2zYkyHVD4WF224wm0T7YbBoz
JNzdn2E3LTZsI+3qSrj/OahCOOMHgD9Iy3PmGQe4tjN7fZrZpr0uAUBROBnj+yTx
2TsQTnUW9/VJaisNkhcsm718W3vAUnQ5sKU2cqIxNXE3MlHmufmcq+Ovb0U19+hc
h7FJYdskIwLeGs8jiGas4w/eIY4pPA3PYONQoFPPO4DUv0P74DcSqSPxxv9Mrowj
dcD8KV/MpgkX1kIJgB2aD4hnspIHUc0b78hMWyqHkfC8sN7rf8pKB9PSov8GTRt0
ULm3hPW1hj83cnf2xQxZVWCJE3r+X76L5uQ01eupZ/PfPmYzxjEYqbw+0KRaL63E
WyX2oN1rqFVDyXcNBDUXjehnoUTv8zj4E3Xw+ltpiCFO+JJEjOWVvMFje42CkHYe
nDJM9WgsMuos0O54WCwosTJhOIiW3YbgRURYwWrp01zDGjn6cArS7Jy8bI5E/Tiy
HOgzTSZJrpxVnUjIo5KpqCt9IFEguqGp4fqwoijdX7M69qMD7czbj8ujzwn+OMAD
S+wNBhNU7ntb6L1lLv4zKXD/2FNDgL503nE6SzFlMv71JqLiQAnpeApWYDnM7eWi
Y90Zap3f8pmyWc64v+suFksyfSU3YQTAZKM0+mQpYA6DQJ55Pu4HxrmnMdbTsEBJ
3Aptbkyksn4rtZZemT4I6DlQA9eoF/aAa9ZVdCzM58B9qspHBsQgaixXq3bvIxeR
DgtlznGKPkRvSJxQmnfNAyBIezyIBOrQBsVYIJCe5nnZWTHtjG+8kSTvoan/OQkd
OBzWoKGx+BU/vmM2rxEmi/tpGVN5AnZnpHRy1h7bO40c+tW08lfcwpscsED2eNG9
UPcGpdxgufQ70ZbZ7ijtf93Dow6PI83KEr8QuzPceuANiaru+6h1ZQhUUTY058p5
WFqyUNDJNOsHh7tjdEGMWYn2mWFk6TVgiJi4R9VBquQJxCjMECVijcHqel36H+4S
FE2518gBrQauoe8zV9rV7gsRWAZZTrNtuMq2U8/12ug9tjdAjaebnMGsFtph9PgX
4ozN6q6atrIdljQG2H/o7Upp8IEwXYm7dVE2/U4e9bSKpWCwVfv/VJ6x3qCdHMys
5OvuytO/qn22XQo5vzuul/d86S8QyASXtd63MPI2oCLrLMtEnLfwJOGT1OFj97xi
rCtY76oMDvA8KU996nCBIVyb0tVvxyZtXAf7siAGOk7L8Dg/1IavK5qNOjm6v1ta
zG9ZWv+Er8Zrnv4yqCUGBoED/WYDiVGBvKBHmKRyeJgPJ5C166OcxrSX1LU//9iX
FqVMC1Ho3WjKriT/5O5Wu1DHUEEeYkekCnB4OMr06Tc54fK1Y9wl0tngSLLvnp+D
F07d9Q6idTHJevIlYvC6y8rPsKbxpv6mxYQidgF8dZfFcFU0+zB2azei2JdZfqng
XJ+KjM1etJJI9pA06fTj6DurpmDi+3CxLiYftbCwRgTBMe+Ov4qPS75Dnmn0LRCy
MPQxAeFrVrl0QcXi+Ux4yZzujiwbjtEB61bmyTW4yQqC42VLnKmmFDd66hqNAnzM
OaIddSmZqEfE2H78nohvPOTAVJiWE30bDfyGsu/J++T+8LLaiJKqgKA0pKlL1XCV
XDXdkfgLmjRCz7L76vjGTw5hz8/KeGl0/WxFD9p+ETU7UCwMbKdGSd1pwd+11GHy
MPVc6vN0VQTvNAeYGlU+GUSurOfmixM/P84VhEJ7Ve0Z2kYuP2Laranu42sqsNpC
VrXpkSBF3tZWLYw0jD7mEJlS1mrUBcnBQwzXbE1he31pV9C8nTn6GVc/jQORlNt5
PGnUZpmot8xPTmirv5bvWDKCpsF9cyYNmbMTGVPq4u7aCoCUDy+PjnoDB8W45I1U
1q6Jo+8P/YpqOXFFu8d521rJwQlTkznQab9pQzAZEbvWw9xMxJIF/r+4lC7KCSjO
thWFVUeVLQNpKGIbOaeWMPhK09YPMk4nvFIykD4m8M4DH5tOPLba1dCNNZ4nYzT0
LVXSnFm3E7DavCPe3+lsRgBTiHV6BkRqbze6f5UW/+2BwFYY9srdjnarWNUvgnaP
N1Sau1hcoHH7iabJRDeDMkIEPPAuIX+m4pLk/R7QTc3ExxDBXFyCeIZKMrbeDjKj
g4hvJT2La7UJ5uolJsaHzeH/FzHGPytffr/jO3rLgCikV0HGmNJVX6954qL9mf+H
o7jNb6Yf0RZz4q8KpaHt65th0I/js+T8vUHXZizOZp3+qothud+zyBsCpzS9IQ/9
rt2cdDl3TFTqpA55+Ipm0T/c12/F476QiOzJ9eis5R9w8afzVZkhEVlfx0UTq9gT
i0KlQ0ntDsIxJ+3N5d7atYjsWS27OR7kb7sZ9/SPUsONVFPchfAvm0WzULLAufj0
Pj0PoYNybDjGRS27aWUMqQ0/IrNFoeMWNc1VdOku/oZfFVZGBYj3pKM/XIuI77Bf
9mFw68j6/F+eb+NTJQ8/COn7X7V+FV83WflnNJhr1tKUhjDWp5OzL9K3xU70vKTw
icDmlHciqUMQb+rgeN3GoTg048kjL8cRs66Z3zAGieKpnAmwyu0VaiZGTIqZL6qD
jAnBLwJkIL+rPc27n8IAe4Zb2L03qd7cQUHzsxFiu7/TR0arQz80YEAyJNwGap5W
TO6fkN+LpXFy7IWyCqumbl825rldO/jXPIWJcTnfzvGqS/h0vC5IRmZAiCtwQLrd
HnyO1+MsF8VyeexbdL6VIPCHmH9QUiWAKH+pSCv8VCqX11GNZdVWrNnpOPw0LFZl
gOojSpTcArR2/kTgP8L6XV3tfa2NtcdLAb1n8LxpBOb1dA0rDdQF1fFlrPOIIYCo
yq6u4ci9zNWYitehEBHP/B9QQDo/Mltg1aQ1n7SwmmEM822BHVYYnRZlEyNNsXij
7a8KSCTFOzQeCnFpt1/ApVXY2eVnjSScExMIQ9lqiBezrLZ6ls+G7VO2fsqJXAXT
dW7AP3KHsorU1HZ35jzsL820e2EDTbBuPL/kK1/XNWqxPCKkUn0C4PXqK75vZb3t
3YLZwmiEShd9Rq+guvcnjAMbkQszTdU8t3i3FwhLc9K9BY4Yz/2L1O4h6gWaRKo/
RrT2xGCLTDm6hrNqlg3MGF/jzokdG0skrPf7SKEo2p0OkD4aMJz0ulbCmOwqpHEo
zQ9Y0yFSdaTFuE2csyd94i1SFK0wiAi/BGYbM2T+8rSAk0XrbjeLGSUdvNZRSIfE
bk+SbQ6HPW7OjH+1TyTap+WicNqIB5x/SCZ7lD9cydwmq3b3MrDERpTWF3i7rUpf
0+2ZATQjWhW2FXE+BJusn0zmRjsW0D5y97rVYNCrR1bfRm8Prg/9qgIemTXC5JxC
JG2+AYQVv/MWDZmPLaNnl3f88DeKUylxFnmQf79RMuTRNoh7UlDKcHBJcalvtpEY
kMPkziCl2S1yKtF7U+tqtyHx7aC5G4eWj4vVt7jKxntxBEwffVDqo7qlRWyjRXVz
R+1ciAh4TG7JESG1FrC2SkCdpncYYy1gfdKfWqL797ovu4xNrKO9/Oo9LCRIctP/
2Nl9iajfJx7Abl+Cf/Nofzex/1P2dRM0O1wEKaKZDJmgPfU3SDWbtYo1w/4L3iEo
3uZIHRGiNjjA4pdHMS1rbvMMPgvMd9jT3ydBZ94UcZPpGPiLzvPVyt6zB/eMs+EJ
95a/oRyvtc6Ch2MJvOdzowjkqXm3beUVcXzNTiWdoSWEHGISsZ6KzfTaXIuQZiZI
MsgX9UpfcjO+0zRsfmSDCuBvLfqaL+aGiWUF2x4aDxIBgOFAYNVH71MJV8nAPBkx
L75t2sgw7kgiusqbttH6FYqWJ+tA2rRAuBLWaMIk0mbYc7+gcGQYWvn2GcOyohGG
QzVXjqgrWb1fS0JlxCiokpNvQYRbyix70MAAkTS7W9taa/UJVntSBmwHT77sF4CJ
dC/BiXc4EwDmX9gZ8hCJuNal0L/9Knq6N11TAD6GjOs6ShTfMMdwlrH7j2URIotY
m1Htu92NAKyTmdlqfxH66a/hdznz2Ng1s+z9dtgLSR8BNtyAcU1RZSfrDiL18Ghy
xf0CXHbaKK29efY+HlWnRQw15y8Z7oi6zkkTpSyQe2V57zAET7cnscNmLArv6T98
qFqqvjSKbL2o0OSui+Bntg/5yGof7PRYqyDLBt6wBulOfiBx3TB1ietvjqBwsVNy
lH7IlrMSk7Myr80Kw+fpWGDG/PKNAoZpT8gn7Exkd9tkO4bx9lS8Atm2WdUdDOdQ
KM3UfW7Qr24KGoT2pk7hk9G5D31HV1ZN0aVTjsFE32KKalr3Ox+HPBudl2nU2oAm
8o5EVGKTheMjVcK7RmxQXwDndj5bgFnE7S55Y7W6aSrwpqqown0jok48YavQJuVf
bPBEntNI260/2TialIFS3vAbKqN8Qmb4g606pzAmLEUD41uzKedYGHu/VGWwQT1F
+RvwqVcILAjAqOHZKDzbzQRlnJzpsBGblo2Dis5xrY6B5GIs6WnjFYCcemxQYLow
AIjgUHNMDhqgkyyn8LjRSADQpNiZ3YG/DdyogrKxhoxtd12rZB7K2m0FEX8w/yla
NW+46wp8FLOUUsHOUgMaQkTxJg1KkFtzNwAFQzbrq6cJqKeRWFML/Zm/HpnmiO3Z
zfeNFB+PgReN3A9JFalFG5xCtSa+9RejozSXzqi/TpRH1mO2PJsXKEnU6cewoQ89
vAaQrxy3zDBUQARP429gtJ5LrAHfZhmGKqa2az5HAsH3+TPUYcd8OkUW9ntOMDIq
R46K9pQcKUc1jP2XvXUAXb9q7Gxk/8+CWc3YdaKhRKghk6WKYTaJqzc23ltXPqWx
+U0OMwLdtfQrfaWw9WjHEn+5aYzkzZ/zFFuAADUKw0sNzVwlY2lykNSLckuAAVpC
SnVoEu8dorNJYl1tq23MmKzk1xN3/lRrc4Gk1cWU0WxP0LWIL6zri5ykVtQdH95t
dOgvKvJ3rSATT9BDFttuOO1qwEjxggLwvAmnyBq/5/uIOVZ6J1JtGRBmUwTO0kax
D6Qm6/swzzYt65D632oZkZJ7lIJqvd1gNcGy9I3xBkOGQYIN2o115sFKvm5duWbG
i8k/c/ewfMNzg79EtyG19zbXrflSMTKXJ+FWFN8iYg/i7L5bjRuQdEaMnfdzwnk5
lIegklUBzSEcoLyEf14zd9m5yKfgs6iQluj/AvIvAWj8SSGajzlDi1JJuEYWf/KS
uV3omM04Emjn/Q2wB51LbVeczh/4za8ElNJusTrX4IYwSQvy9osttiqlXlqioaoB
GEcyH8yHSYm9bc0Zf20lqhbmFMvrifmW0lcpogT11OmN3H98dKnqWuasqxIwbnf+
UIq7aYAekqKsqvYyrjz4CDx/XwqVCGCfgtzao1ZBxszh1Q5Z+2JqJcVvPxAO9sce
PogTRdta7IaoHR5urxdjUJNTuNRiyonTOSHo+/I+4daTIO/+4aJ8Rwu7drIW6ImS
6O9vMp2RIcSQDIKQazDHdFvtTrJlbs4ooJHF+yEHWPwB/X9KvaecGP8DQ5nZOxDn
6JUrJ1/8+8c2COJ4R2x7CpjwTc/LCR0v11gwCjVzHl/qsR/8PElLMh7w5Au42vMc
lCIeDIWz+Yi7FFJ+v1q5LabMWuRDS4adsnMk/yKg7WyVJxa1/zipmL6sKvWdzXFb
xhjbyzpL4tODTow7BEdTqGJEs7DBRfbRIe5XQ3kmGxqPgsMLYvO45JeRgtuiCucI
lRoltc/dWZDmc1HtAOUuFkMlx/ijd6ywSt7tQZC+CbWkcS9U1OTq0r8GpD05jh6n
YXmrhVSRciShsQkkIMwt8qUfzDsC839zBaUGSlLhvIal4ZA871Ycsd2iwMBdAypo
ISKojN8ZHLMUGbI6ROz2Y1yF4dY3ZC613tDKHrWdE0Y5SnRRnIh0Zrdqb16gzABG
dZ2Sa7RHoCSvj1rWlNHEKb9d09n3ZIwhlaTJcNxKy8iXItah7W4ZOydj/TAYUIeS
uStFQx1IhAsyHlpSOi9LPJrqrybq5P4cV22y28yy99yQSU31YVbsu8wuOEjUMy4H
PEt+k0V4MyJeT9yr2LLTTJWGgxc1hxxrcY0AfLo3A16FZA4cCb3RduhBEHEjlqQz
0eHrmf0zsMEeYlLZn3vAMVsE7YcNEm/6bYPyLlRu8/2hCJ/vmW/mMR0yHUvEvnAj
08tyiTX8EbZA3ohF1/HmCbxNiLOzWxDu0aAl15PRUBSk9c4CvOYRRoPEbkjBd3P6
HcvU3/PLtXNCtfMGfy41l6Cst5CLjdr2aUOOljC5J1gxz/xweDSJ9jUCl3wS00AA
DkayKqjO+W3dMoDFCFR3hiaRv9w7PMf+MbM97/OA+2PiQp/x90KopKhw/+T8E5Vf
fTBnW0NAZJrDCYXJRwRbPnmHEg680jwYs8V6/byEZzg4LmISRbGOJ3G9Dxf7iPps
jICoo/VNT7pEFJHUM53+7maFyOWfc35kmAntba3fc2mPgyclxGalKhRUMI1fTvkz
2wsuhTFeXPN4D9b4sKVanFgt+iKA1zVE69K7b1Nbgow/IYmzh/pC/22ROFE7/AZk
/SpPm2v/9NewfaAOtQhevS9h/MPRTFaA31TZZxUhJEXSayABO6dgHpVtoMAyvEZg
axl8AgEOhSGzgbkGCbNmGvO/KvhlJ41xfoy+q+s7QrZLVGZsgPnX9yKlWCelZmE5
7gR6HHDVHOa0dC2RZHEGMWYrtQp9HZPT+jAermPqLIckECmoCEllf2xrChhYyqC2
0uubX2OpQJ1nCtimvEg+fiBxdyKDK5UQjc7wrBfAGKkg8GFNTyCyw2gJ7lCgiT8c
OK5ZEY6PFqb8PqarsAOiGIDepxbEZJxVDZNZ1613jWwYEPcP+IVyKLmOMb6IU2lj
Taubn7pUcHS90B/lv95DOYXkF5WWONI70dNhkXmAGmYdmCS1VWQqSQUnymT7Tr23
GZM+foLOJ0D/5z2kt7K9r0VQYaF4Zj0hXzRXZUB3C4pkKV8jbDkzmjDgYizpKpg9
nUTEGuQfiuzvVIdhI5GI3bfN5dxlUMsxISwUaxKI1GDoJwQ3RJJukjKu5ByI73gd
F1VPjnWmwoUUi7eo8AyaJdtUyar32NMizI7Jlc5haKsAgQL348pU4jJ5bZRiRGXM
kZxUz/HhFzYdRDBvM1hBIuYiqs9RQyIFp/T+lqfzEGlKWnb9zUHVRsrk350bLofl
41n9E/014XskIzMEFPQitTP9THMwHQhb3JikPk3JN+iETnZpf0TRL632v8rzWFVY
8ivbau3C36MCyy173BJtgF8TrdrCqd5yd+OIHl64B5dfZXRXnJWSAKgahBqnW7aO
fFsmAi2gMUU9T2dxAN6N/th/ufG2Z+aqU2oFpCb32FF0YLEoJDVIPKuotX2G8dmY
+OYlThyieMddbGB+TtC0RslfQ3Jb2De+v5gJAyXTrQXmmE2I6Z4ZqRavyaXUL8W5
jWeC98UEQ5ZlB/YgaHFwOinq1ktyY34SL0p4gfBrGMOjfq5EfoBb4XeiC2tsnKbk
9vGbrPxY4uvtQ3rWQmorMyDgPYcG0yGMSWR7YAJjZsWrA4ZeoysEFiormKOP8prP
4Mq6gq3SqgjWVc9daA5zvhTFc3Zv7c6an1vK8pIfQDphAVtloOxfaQvMsUPtAUkT
RPNIkeCrVSQwU2d3eweylaf5RPwTCBPB712iMYwrmhz64dPW+K6CkpSkOd4EBezZ
C8F79Xh5YAGvHzhNwmgbTb5Ud+/6fOXfMYKpoYGQmzXhRB+AvyoW3tI0wH36lZMT
U8thuGRRXr0b42Shj1QmSH9QxWMTaTdsUbKAGTIyY8B/caCV7yYgH6+tZVtJYG8k
yyQ+jZkG3ljxTUJKlRJrsNfysJUjoLDsXy8ANoGfkLqGfy6x6rSWzoyyF4Ec8XEG
xGsIqNfWgxkK4p1/ThBaiivMU27381BVpZcQ4A7xxm9+3ef3IxCtQONEnbggld9Q
lfbIdUVO1tcgxpeUHMi3VoNMsPmpoRtgL6HIidt+isb6y/iG3OCVC+P2YZdl0sDH
tCcXcIAUf2is44tM3pQwN29sPoZ5pmM0AviiZs+NdJ1qLRSw+mGmOA4GnFGRQsjM
iXQZHAkYYkP596Q1cPXM71Cb4VvPj4lqgJ699494dLU0q/8iJ3lV4RlF7tQscI2O
9LL511W87Bgn/uYS6rSQHAfO1LgNLPraP0e95/rIquBYDTWJMvFhQf4IuAjeD1MM
bZ5c1dzNAVeUAl1n3+ZEfDFSa0EvoKmmyiaSDRAmsX69UmwXyc4ICI3fdVME3x/7
uj71Re/zh5ycSrQwDZasF+nlJguV3kLhCIaDH/FJaE1lj0sjg6PVL4Y4dNXr+FQz
sGkAfcWgeRfkHUESotDMg3IFVgNmivJaGjdK65aSFVmL4gWYRPPaj4KdK/7hqJr7
8oEgahvP6D05ofxKniAvu0SEzOMYSlSfRTKk3g3FS5CReKGtziuvrGeUOntvkSuy
uEeOn+h/rO+0W9fFNDS61X1PbilavWjQ1QDaG/VcXymkx3rNi2Z6S7reKUMQ0t5Y
MaMOPPk0G8UKuTDvO8tVDf30VymoZuJX7v5G8Z1rwXwEoberySpd3wR4jVHAIBcH
07FyjXmDCNO2ShOCCndKZ/VFfC4sN6w9262/1xXAORwaQsPTMeD8ZrcmrxxZrkIw
3UvLqnOTsQzaojP3GqRhdN21Lsiu8wqhy/o/RYNALtUDJWTTy/WOFMEo/OpY5RoF
RYwruKLUrAhkoZ6jyIsGFCwzNbBfnsQ6Q/jcJO5MYMLGo3qxQIFaRlwAoxxvSq6A
AWrTDpaP7B4GphrBW7xt+t2cj6vFsXefCNYJOMpTGSmlKN4EhbRUZYUS7q11lMUD
S5TeaXw4QeMZqpXV/XI0BujmxHQrgL9rEVC6UtNblNl/meIBDYKbg8l/AM607b5F
E4hA8Cz5eZYfKNBfQ+5XliYprhbD/02qCMNls674bWThl4eKyOi7qVOwcUJygNoW
DQK3bfCR3ADvsE13ves5ma+iSGGyooSPHCxXIUsXda7GTB6f9VWOH41WQAdwowpc
flrsPFcIBwegp+VR3oWmPOpeRtHfWblZjmCMv1weOkMqBQfrSwFr6slRZl7er2WG
djJCNaOzcJ11NDQZPRm4M6ybgjVQNdka3Kmn+gIqGiC6Uo7b0dAe5ixXolT69EZX
iyr1uzSuH95eQOIG3jC2ON0DzDGAvgM4z7o4NL33BeAVDVIfBVBPUgiN65iOP/+/
9vXKxffoaVkCVD8NoELGqHi6/FVuwabooxRr2G2ruJwvpMSdRSBoIz3tLpgbsmBQ
/8z2QFO2eWR/1CAucllC3LAiDjc/zUIT9zOlrsIrIdfrjNgOs8XxQDhSjPZcON/h
1WJXtGLgI5MjOSBuvUGIkDzh48pBRxkvHy5+jBhl9d/Hd/em/N+9/6xnVrCfeJJP
2wBTsCDw0v36n+pxLgnZMCDIBNJj4LIOdac990xfQ43RDeY3mI5XgRZCyBnXrRuG
kTnXwwhdgm7Xvuhh+TUHTeQ3/fh8DsUDAkswkF9kwqWpsZ9zX+PlRchs3XrV0tYk
d3QQPicT5hUYqtlDZ5OONfZdUOthWn1tG0noQSrFYWEFMGGSxfohMxdcSUcNzusx
a7HJv9ofUr8535mytyxOF55ZRl7tZYBPRSaibmWsz3wBN5AvfgHPtiafZ7r9hJ3I
3E2VWBJIe9YF+W76QLzjkr4ZrSZn1SjWaeggHdTPG9SOvZoS3MGyHnC9LPmDfhd8
wGZpDS2pznvyeDH/+B8zQHAv1azCL30JlR5MCRqgndiXBVaWSCko288ddEvZJE3U
jnOmaPZPQXMPFOHwssudky0xegSXV8r2sNGo/YEOyBnAnuZFvddOg411x2o0sXlG
wi885uobybXtsPIG0yTbdulapbH1V+yuhPTwxWT2lmrTtLrhaS8Wv8Gsaq7iP1TU
qChCqgZFxchiZbxmZyN6emY0SZFlCXxdzrOWoZc1HF7g/de5RNJWdE+AOHQ+3hw0
jyN9MSDtKOm+pC0wMiVbbxEpEop+cT64SYHmQ1nluWnS40hGmkqNZHiAumAXkgZB
iE7QSZBuz1BAUuurRyr7xOYT6AZpsvuw8KRmZenazYpjvho/7UguNA88RQopeKHI
FhyxgUR299as0pOcbJqoCw8tQrVqDC5GavcrpWDs4rKMpjbZXrpTs0v80ueHJPuY
MuTCAbR+wg78M6hbGiWkOFiMM9NFNqZXE16H6+jub0QRCQyCo9u/27TAKwx3tayx
s5pV7+meSsBTmeDakNsXJgYJUrJspChT/zLfd8Y9CYy8qCXAj3x0SbSo5xyiY4mO
eWYd2H9sRmMHJY/ZHPjr6ty7GgXHPLvFwM83PZnWVHh8GSEIYYbHSaPal0JRzhV7
3NCDx51i28jJy4K0RUl8yIOUjlYYTRygd+FkGhTw5Ur6jtbSFVhZxKqMta9+zpWs
rI0GnGfOQdtIxZp1OP5oZ8JlBmxfihaaQHqHsOjtXNqqiNIKewoS5JJv5LTQHSM8
rZM6Pq9Zuh/MGS2tPmLV2jSb4/lN0ORr9GA05HCHtRTg2mfqHlsqwl0s/QLPAAzP
uf7Vw/XnLotoVP/NHGFrmVGMAmVYnzWJ7IJvwCywrxiI7ff1s29hUxdMsqBM3lmr
Dz7ppSiUOA/koXYfQ9X8tIDzCR8t42sgAnN+pVfau6CFSYRYH883j67EJ3vvhnSA
drmnzYYtDLvXBrty5uWTtxPHd51qrhKgbUk3A9Fxxc+EHytIsJmyF17QnbRnymiP
qFo5mIoVS5qdGu/edOX5IwZpKUrIpD46V5t3mAdHmFqS+f7lrLIw35ox6WQcXRIP
iw3u/kX8sNVk8KEUs+fomzcv1SPglVDczLJr3Ojv4a6fpFdrDShSKLIo8kjAwQHM
rcDgTr+QyDM9ieT05/yiFeu9BtEDuxVCZ/yq2SyVvv1NtWUyX9gCjHfSbOmzN1RD
2YSd/VLdNJGqLObWdkaROPEUtjqJLa976uzuNTT5Sfa3n43xHTrg94sdckeyHWy1
/EVeRB+Bs+sgflPHhjAdT+R1RdqJ0NlEa8qZQeIR5IjVbuMm0A7BLaLNIbWtFFhO
+VeTRxsuJ1eSWkwR1ro4LFjcbpwT84QOyKHY14J7Q4oxdISQpbbY/6CAwyHM62OL
w79nhVSV0tyxuoG9Yr4BGuTusWiCofvoZmHPGeexA1Z+xvOPjyqlkQNDotiARmxK
+wMl1T9wG7dG+z/X+Gzr7noVu5wecXrNXYKOwAMccxU46xLl/b3Gux9NNXaCIzpf
oLnhfziHarlRL3PyLw+RrXWUXHteU8rk3qymDm+DAd5GYCzXPqFVI515rqMoGUel
LygmcXkLLEFrhBPdesQZknbnV0/fAKaG+aEREXCCMXj7uB4u9XiHxWu1fVzx3VW8
cZJZAPPwbL6IDaXuYqbN1M0wGELc//UtaDzIar+UFWZIiwmZmSX5kWRHK+oc2cBa
1Nw9Yzw5+J7zJC2nqgSAFkjvC8H8AzPOhQDYP7woiB93O0M0crVxlfR5cOlUOpys
LxPeObZsZ0aY/QfY0kgVqaWqQi03CI8/4m51wvTbYDLEs8RY3hZeW9/ys9vvNfUx
1bz7ZpmYlMWDCEa8anLAj48FLlILrg4IxsiDNlkrnoaMnUy1WZurKdAu5kpyGMMy
81ykSnmeSRX6Ggp+vQUTrBW4d68rONyjE9mXUXDELZQsaQ7UNiX9nV9qJhO73RBl
n5MwHYVThWjxv+w8QbuRf+SEQFjloorIN2VxlCtFejwHp2CrGzfZPM0471SXwlpQ
T0GOwm9J4WEyBCwPoylSUJrPyl6d9a4L0nddcyqARsQsfW7iWM4eTPgJCK4TU1dI
Xt8POAg/SLnF5+yDCKmii4jIn8XAkZ20sF3J02ipQWTpYCDY5+kNo9IpWNVx6Psp
9/xyjAf/Ns1yeD8J/XacnBcoVpMRaBN15twuM6h3/GWleYZI9dk/6V55V5Twd37h
gfNw7M4cMWrdq+peDi9/7rGOZIlpWoIWI5ERZcmF30ViXyE8mBSFbTi32FmG0Phc
5tnUqTKuPlDEhqA+/Ed8g1aLg/YL95LPZ7neqyd3mf0wNJcNpuuIlq1qS4MZVKrv
M+OzJdr+fpcDuziTAqax4dig4zljO/Xkfr84fR4m8bdNI8/rrLODxETFjkmTGtYC
d6hwTPECU23wRSnmA+l8ELfmWqswPNlNYESOvtAmmzyZi5CAfRv+QelWT04zmXwj
QKTNkYCLUWxWe9oBglnuAQlbhWMHTR686XzdcpZh9KGI57Yf2FtUBir/Hkq85mYy
Zv9YV/rDGC7vM+KRF3vtP7OP2fctiw8RvTd7DH/jukZImPbS/b8i2sCxYiMc79sZ
a885cXLRQnSkwMRuSvxugRUB/UbP5LrjYNwW2a2LFhKqJR8dgv9k2Rja55oe0o33
hr3Hd0xhsWW4/TycOKuNAthJ41BDYQniWzUeBFqQJlIdctD/uGVvrN8JhOe3U7kA
Yy0IdhQL52klR37J2F74KezRu4PlC8fIoLcxPqVtQJ01A0tMTOiORwl0tG5FN/Qj
Wt+ZKo5TGZUZvntcquNe4v6NZgsXe7ySzYIe56kTGpXCSXMuC9Khf6o01dqZzkVn
4g+iVwmv0sWKsh0zVzZ8jyjTDoNsoI+Dk8OGo+9b5SO78bWSOGx9pKbrIvHEuX16
vn3JFEBy0+bICqbMDhCcoZFcKoCHHw/9LhMM6grVIIoW/lj7aIpv+mKgG/u0IHvy
G3JYuXvZeA/Ffaud6EaE64zEkGCnHNgNEkUEpR4RJ9+I5N9x9pMi5rBWR6hIXhz2
NoJn8jKMS5efqfXute6g71hnughr7wwbEnQfPzhSJKYwAQEQ5O7Y1qb7t7HzjaDP
t7GzUxgi8f/vFFVLi5hqixMbr3p3gtKQBkGUdJpmAKdqkDA+jKACnRXcSaBlqpkN
bJMwEo1eEVElCz09ExjvFMOrAZP6WEHgyJ5/4zWASB+0InHnU7DPIl5yO9oGJ7eg
TJ4IyQa02z2EtDX4OOVUHo0ZXgWKWLXzhPLNm+qaFjeNc6+MWRpdu8cGIpiRjla8
wJOn6xa6d5esTRZ1XYvmQAAIvaRIJgelXzvUS21J6dBSMLaJdt480wr8v4dIXmlP
LV+uf/I6RN0On010doabFETAX249cQhzbA5u27apmvVKPCycjC/Ucw4/Pe3Fx3oL
irlxYRCU/YxS52/W750tZM8Zg+RLxgo2FQSAiSsfPOOSfRkxLL6HixoDgSFe9Un+
iDwl1mwn8jAebs+/BFgbjxM/p8VZfiY0FWF1B0m6psfJvju8s2nNOkC9zf27L0ib
HFd2zfSN0mA4J78AqOvWA6Pth2VB/nU7T8Tpc891MuP2swF8O6h5bSho28mwxyWN
zkuju2gMgOtLHebPdmUVYgAO9qz6VcMebS4CyyGqVpoFOo1muMOmEP8E/b25htUh
Dm8gXVwNAyCXE/Avat+4YjCepZvd3j9TSqSrGPS6Kw74xauUEBqcNQ9MUU/xFbjD
nAkU+boOR5y3wJ6EHDka3tIT/9rkjZrxrIddxmSRqGLO0ZVTgGZ59TjiCOeYkztk
lHelbYv32GzjgDdpIso1NuYqMuNB6gp1MlY7S0yu4llYGVBaCmnw5GFT72de8xxA
f9MnSvnPdem7vMs4SxapxZsRL+3Mb+MvEiuGN9kCY2Iwoec4g0zfQxw9bjyYsaCl
kU/x34ltJQeVM2+uH5l4ON9Pgvp+wf9gAPH+Yh5MPX7UinJdnCkh7NTP+PBNr8Gy
oCqwVLkDpTpbTnPxkxAfjyB3PSqF4/+f2DRfqEldhBDaUKjuu3SzAng9wV3Al6qg
wYJDGLa814TxVGSajB2EkVjDUAx33Ye+L63YArn9lB0uSwgUO5KABE0qdU53aBVK
rpDTh7DDw+UX6EqNJTke+AA2tcB3iQyXAXkdvmSM5meq4wjkbqVRmbsOvM3Kgi7P
kgc5D+b2YAzaQpQZKJEKQzmqRAVFa7N3OJqlAwpV/C+l62TWYSVF8mzzCuGFip+3
yV/UzsVU0GDoR23WgFAFmBXl623drgpo5EZLU3vrWK6qkok91sIOSRMLjS5+0IpX
mYWzpZ123xdeLqpjGjuRO5Qmm0ECWBQws3J0Jdz0qE976E8U7AVlx9P2LXEU0OBs
fULPayYGzDPfAQeR6UGhnsjyTRlMVf6opEKSCzz9AfAUA0PjxC1kIqZUAwLJJkGO
wYALYZh+7t0ZYm3lSKO+GdI6a+MwPIJ2wZJrxtJICEIwhGvQkq78svCzA4/W37y5
UURaDyV+IAz+50YWnNLfX56MHyvRxFXo8gIkc/RQ5b2W+4LCQBhEuM0wjY8bhq0W
zZvtbRRM4VpULtfhdPat0LarTkfhuw1il/CxO64VtXgIqOpV4OS9+OoI5jwlRxXu
tzQdhhivmaUEHRs3Ub1fDXNmnrcmlF34y0o5HzimTiu6zhhePfn3cRvuMu/Kn5uj
J5LvObuiy3Il/77z4tCTUB7Ri2Owlyv2fdgBAjQ5QnoZFJ8Yl3cGONwC4hTFwZ58
pf80BUEvVoG5g8TJMX2ig6XMOnzN7EX0JAvB0FxPWiA4Y8YNlzMa8F3lV1Pg1Dj2
32rbQNZ5fMTuJEroiSzpV26j56c26WSzt/N6WbXy+ocsd91kF8TIFe4HkL2DyLYC
ar/7YfGHvrf1eSZhjiEWps+dB8oRprlqt79efWiokKN2QEjCCQfkVXFPZRXET3Gy
iNZylHcaY+ytL46zCtWeD736aUkdqdKXv1pUOKrM1K5EB1D9od2JEbqaBNR7TQ19
NsN0SwHGzW6Jq5USRY+pcDLbDsq2lsMWUCh+DBsVHFDz3QQj/eBBcUmVSdjqD1jc
uI5J5XDw80YyeCD4YkNOARPvFxC5wOkGRBDOV5R8INcCyvX4aUjApWjLYPr2kNnt
JjIzw4ah7qJ7z8u6kFIcqbQdgPewAhvwmMWnCBGHyLDABCE4FrQwm4kCovqnu1g8
w58cLiHdkRSGhjwF2IhDpVz/sH0f+IwtRHimvxhiapVgXqVZjQkLKIphmN2Rky/0
I6z9J5iqmejNrrWhc6VgliAEUkrQWEd9sBMYOEhPPYtXRr6Kyo22iAbmpcolSv0N
2NzYrWrnZ+RNgr2FrcAuyj5mcXSkqz2YKjMwmCwmJUK/ETg01b21BF8Kl3ATPVRd
qGDs0uI95EhsmT5eyN5d9ickWr3afAhDFnA11NLc1h/Hxbs3UFNOMzDWQ91BjBdl
0thVJkp02NrjtV1L/O4K2d2Hq5p54GMV8SEpOiC5+B8X6ZQlz8/m1nHIlP23Hfwb
fz5P38rPUEREC5YfSBvpS+A/g+CcctMsT12JrxqFTPjJpBEfVWIg82Gr8C1S+f8t
8OBVzN7k2ahn1irkxiOWx1Mcdcg0DmofxmwLFhrqJ3ZlcyqLaGJBTwVZKtyVld2N
mjRKC1a+vJ2siqovSYUvrep5H2TI69wmCoOeJhjKplXQSpCbNadLIGtGT8FeOm8C
yMpDWDgPLsA56TWSKCWNrpqwBHBNqkDR7VrgGW4yw9IsMbIh3p9iM6HuAZmvMnlA
40G4veK7w40CsEcVOEUdtWqzVXTJt3ZYVxlrDLSFXAcmYmgOhgy/SRrPVC5tISC2
SK3v8mATTcayz9Yf0F1+Xv680QAHuNl9eZyoBT41vKOtIgsyMObv1MOxWWqRzXq5
F4A1I6eJwz49eF8uNmH9fLU2RBIvpsxCfiDWsXdhrBM5UD7FQhuDRRuTIjukIyrS
vSV8EAQ0F+larr4SlyR9AUdwVtBR1Vb2qLtY4U05/CNBqAec976TKLCUKgj/PjaM
HFipeQr0WWTOoX3+7IQa7uyWi3FPBh6710vbHoU/Kuc8iIUMRIvvoYU74QZGtBek
qE3JEcKKTW04EEGm3a7SfIiYu3E9oO5DstOA96CSjAPc879pHN+skqr0iOUyMZJt
3Pz0W3Lrp2WzavXxTU2OpCOVE3V53S4vtsdlnUeyh3Vl1qsztAcpLnODPJpVAJgm
ZgxjRUT8nWlCU0ltawkIaiGKiJZhz3su/HEQ26LXAm9IIMav5UGM/UD23GP4rKIw
4z9YhPttBvSSPkb5JYERY0p3sfBe3xrb2lDn10jX0rOy8Pw7PSQr6HQGlSrM1GT8
rg6JqdoYVrVBUuTESZruN0YISyVSG8KibhpBvWUKHXF2ECYIuO88NqJIngVsqAFv
rHyTnIDlrnGnf9ITMXB0bOA/RFK+6hQrMRB8n7CZZEfKTjD+B4tSRb4t3988JgLt
ZVUjqD98XahR7V9RDxBuXnuDg5tXvOpLN4GndNB8RXvRPhRVwNYGSP7pPraZLAav
1CQMVanEV5HkWUEnADntpBwIPVc4mpJ3mSmCw++8R83SsbgfMj5yZ5lp8msAKIJx
aJE3foQsO77dP8mFrQn6Zqn3RH6f7DKBFKXb6kh5X5L8yHxkgaywdztzu0z2dN/4
5Ghm9DG8k6rnkSe12q1xHCsQYao3cHMDi0ye21C116h/+cMo67TB8wACRL5QoEzP
q9xaSAq/F942OSazXrXvAWgooFzZ29NqHs38aJIfp3paR9A/COhGjEL67EXOJpOv
CA9pSnzYhUND2GsR5s2TZEdgB8TQXIgsrXQ8GEBoPjQJruKjX0Z+C7M7YztRNCsv
98q52fOfE+uhz/Zt7UzZE/pKxKUx04XeWkLPY2GTHQukpz+YfVjyFdn6pQcMv/qR
7ZWBUrp/9kMMdukBw9+TZhoD0KcTSOlxQevBXxcWwmu/v1ioJeum4BbpbGNZhPMw
AUqE2ErvaGTd0lcsmHg9KM6mBDHqTiVXSF2zsjZnlC5fYaI/kaGPflS1wtpnr9pK
ChKKDBqlSl4rtwkapkX51LNbo82T/r3AhQCEtSPhpp1jLcej2pKDs3k5E0YV69My
ocAl0IjxdwGkc9Mxc1FugD00O/y6we+crjwQVePNsmvlhb4ZbcKsY15lTJ1SkfTl
AM8aVSfMMMv6Zlvo6EbQd3qBNOiLFfs0VUf8hCE1i5zjiy67v3By9/aipkwBR/8E
q1YPS7GbYqi1HZtHRdrAbMX5mFrUWjydZQlqf41owaSs3nzDYU5rBc54BZcVBh1d
8zt0eKNsUwEwNIAm3TvX/GyK46uSBDPYkeya7+IY8SAWSsgH6kDO6/8U9IMQbMlp
KjFR6eklP852Tztxqd9XiNJHfZmesMlm6RWPh8gwrScpnlvYUwjGerU59h8IVaPY
Lzq8JGEndkwuCkT4Si3Wxb5YRZHQghrshJJBvbELBd975QfK1WJQawrVtao634qD
/2OR4HfB58NcweIdWsN5+tPnyGwxYmat3q8U3iGSz6R4d916SsBr26oAHKtI+hVU
+WeSUK71VFLjauDdZ0tDZIG7nHxRqj99Qy1odX/5E8Y+FnI/f4Az7XzqjlI+gUSk
bdGAKtYvOFLW0S2JfD5yJNTJdc8LUFYOifL9Fgu+M9cW9s/gHi9oTN16HCKd1cHT
c/+o7f0r3oZrJmo4DH3IEfQ4SUMwRBEipk0xbEu4+pKyuPFqrmvo89QjzM/wdROf
uEBAvcgrktyWCuhvwQeHL//1rlXPPcgRFeWwi9vxUxgmsmVBiHtt9BVHH++WGAJT
Oh1KrpdDrxN+9OaFF4ag3t708F5agOvLkEUnycLnIlQWLmqT/bXoNmaqGOYhWWUI
9OT/1ScvZxQIsSF9gPUFKcagSpxr5PTvueED1ARrFBqXH1Obl2XeRZJQOLab8U94
jiWveQzdb7eD3zNZnPKL5g2HCjNI2W4JO3VSl/wXfLcg/eZEB+FMDyrb50w2IlMg
BIZ1103fRiEPsD0i6qY/AaPRX0sTCbSn5gFb4WUU1vUH4vgynzHjJZzESgFjMJFp
b1YnMZy0esWHJggZzKaKPCgP7pUodViSt5TVPjhTlfv/DkmSqiAVOCklht36YtLm
hgC/s2IQ9IuS5kbZHLaxGQjmjgQ366O/1qgSj2ZYOV1heX4H9v9apuW3nRamLBS/
sP495SabN3/46ZiZG834n0TiW1Iqx7RyAdqcMYcAGOrNMV6ghGsYSxkHoSYYZVPo
xR0eCzHRboD67zJhsOIGkFM8WEZMHuVXce6+ByzMzV1EucGpBZhPyjf5llmtfBF+
DZuwbTDn2fAK1kFumTfSZB/1FnUM4zV103hC3MssHBgRg4ENno1Y0Mtn8AOyj3QS
KcyjOUyCn2VifgxfUeJ04Dt9YkzK9vWyTP+SDmxZml/ojXDyoy7eoA+NURji5pGw
wvY1AaCR1RFnLxj3i7uXP5kGkcEe19EcR/dXDklVkEYZKzXAB4ssIQzMLmfGhdD5
DNyk47p7QskHQAnwT730Yk6Kv3aJcbuiHMXfoP+nB7c+33dWAOiwkwNH5UeSfzgc
Q9hSULcvohRKCCoF8r010WOmeufL5xtTfbve57JnwwUerGbjpu7FSaMSn3dCBWk2
HRyK2/ODmv3DQz11O6vtpOwX2Div590UK6e9hH+J+2SIhAq3wztohFo2VYjTeFwg
53p9X67sxaeFvPxDP4KRzHEUHkXRNCCGSOMu9fPZ4YBOsbdZSe8NCkf75k4AGPKO
TpTp2NjeSARmhSl3WyxwcjIsaaqlicA2kBHA1cQX/k6JeVCwSxwp9eYqYFzyFc8+
13A7qJdX3A0AmWFyuuKdH8J0eKwNvqbHGXhTgz9y8sI3zKoj70iZrdPy7oeUVJJU
p/8fOchLNJ22C2/L2R87Lr7zGGwN5pyAKPFmzPb3N3pEQuAiGm7y/d9viix6mJI+
TsHEiqVCwB3P0Ilh1V2bmsU1GoBPd34msXpdbaUNmk6LBP0LOF2Yip21dt7lwROF
pHqXUoTSci5UqiWhgnXFA27mltho+0+plZTxAELsw6pfA2zLiQjuWWajufc/jjM7
J2wPWU2SiWNaXolUNYzxQZjCc6RqzvVYQDR/hXVNRX0m0b8rjGPg35XkVX5XFzAR
KYcBz+ZWvpB9mAmGEggCyjXsIABv1wREaKQtyUdLqjOzLJCR/9Oh1GaFFL3fs/pq
v7yKKyG7NTbhOiuicAGJ5stNmehKqohSb10/v+qNL+6nPXm8i0uRlMIhXvBiXdXw
s8RrCXpqrEapl9IvMSzJV+VQfnPTpBj5VzIlBa9NzhO2vKvYrVbJMVEu7MXxrCvY
HgyX9yclTcT4qFSUEeDsOTtAEjNMOkkJtvzOVJ9jvAxDhYCZy05Tt+KO1FfEOUt7
QGfiozDecWFlvFBEsOvMKh5EKoeBy1QDqWWdWGNfzdMbyUZxKByO5fTuoCzN7L0x
mc99ERK2vvulucLz64a8FJQ5Y8MYjXrFfe9s3mKk8OW6boeVZH42kVQHztCha2KS
cd0yDh6M+rbeV7NZDiULYiRNhIBTNeVl+IOt+Xs+mpV80FwfPLeryU+wNSoeoiNS
Ant+SVfRZNgmtEHX8p+MLbN7mGdCQZ4Vye7/WdUlA+11PSRVXeIWGWeVU5Z+I2GE
UtnJtSTbe2SjKZweHNk7K0BWFAjBNobw2pPbJdTQXsoQKRhDfCC8Hbf08YIfYQKO
qotJ7jjRVtI4UcOqiVMzG9rR52mtV0aamLvGiCL4i/xeI0JfxITBoCdk6HX7K2bg
GqdNOrven6lme5p8PXST6594S315KDRSCN+Rd0KckX9ORJIbRgNGX8YdEvTXW6Aj
J9cIAp6OJ5pQBe7FOIdyuST84bOjtaHTaQW1KK7DqRHAjATCi6w7Z2g0a/Y69c2/
2cWCu/DBdN5VL+ltBo++6Bxeqs2o0xoyusDtf8LPFRLPPh71PwG/ZOFzEqYrixBD
HbLrxXlq2ghfRPU5Z6i/xZbo3rNFLRCt2syhPiWDaT3ciGqBNzKgK5wn5uWqbGYe
EOV0frYlbBWvc+mXDGm5+5IcA7VEY3jfBQvSGjtrpNhCRPvAhDb64JPJM7zMMzaT
UX9bXxASLiW5AvSppOZ8n0qLDzop9j6VVC6UwQjUySlIFdP/onAN5HhaDHO8Jwaf
TX4GLyrbQckagcsQL/mDbzuq0NVUJtXPUedDxqwp5g5GbkOR9/8S+vnfOWkWaEty
LYpv0/T9mxVSTrkllXzWpNrBrXfuhVGMn6rtMyB9SKIsyfReXBe5Gy60ZrX1Kdfu
ddV+FTNTrQAGvwI50Bh1i2Bo4RppHeRbBcmh25dAR5OrEQkJ4OXG0MbksKX6xHNt
boaJGFW38+nmuNbPcLYqIuAi5ifTu+iWGDhYKTxYexKfWGB7gpKD0Nor56ZdBlO6
N6Hnpu3leYwExSjaarPfUGzvdmOg//PxN/XsXZqaB9cudcXCDxMBqB+4CoIXQBuT
h6GLOtRTfv9Zf4/xzYjSkOo6OFDEEkuz9ekqWYsHXX5/YULWcmN0wSDExi9y5NBE
Xk3uq+QkO03cDu/5pSdJg+5toKhhFEKg4mQ5FSCCibmIZ9c9qvZmYpOAPrliHJDL
wtlEdz//SUOVWZeCKRTw2h64hL98DWAvJB2vdU2V0izS8X7sg25YLMKm3uBHdohP
zczFsezdp6BpildCsNaKv1WpLGudNnYSG2XgNC+tupRKP+87Q49MrDrHtKaGZbIv
ziPRiZjV/27qJzBRkDzqEYLjyNnDPg6DlQ5AdQ4rYLc2HpOzcRGV2a0QuiquL3UO
gU5HGQ0LXcwTw2+Wz/y3G6RcwkZFB3APZS3LRs3/y09sC6J/XVnxzMRavFnW8OMa
Um2WW1ekaM7XHYow9sIfLXIEHKicWXAlzUQDaZsSRS6uq1B32MrM/3Ia8xp+uZ+G
Cv44s37KE4LkYHn5CVUFg9Xik4X030haXkjFs6lNdNsAcloaxZIP/7VK1Ag4+wMu
aGWkpFBMjAlPdXZmVH3OmA8KvBwd69jPBMvb3FRp8QwNoEE3w47MCtTA5h9EKkVp
R/UyffhsNpmMKhjV9jwezrXFxZqFnWKXv+ftMPPQPIOKykqfYv2epZiMrCa/jGyP
DYI8SEYGrZdPFncmgLHWELmHORI5bjAFj6Aa2W+07B0PYFTF+NvhrxpuVihLQu3D
AACHsSSvklYfbQBWSOkWeYfulSPJKzcx7GG40kYM87XHPQoTxHgW6nL1agmT68hA
F7Oc117K0l1/S1HVFjWdfxPu+4IH/7sOTSOcZgwX91MsKO7A1ZxTPa8lx41Y91/M
4MKHemPPunB6JWR2yJOQsN+jwG0Sl9dGrdixfIVMdsLyfF/A7T3sWuuOAIcKkvmm
7xXXPM8o/weR0EqZJkYAl5QCj95EXl6iJ+N83wWjwOpeKP1nj+YMsuWDHVWTSWIC
BV6Jyfmzjy9S/zQQenlUobL2T5+D3t9fEUjnl3pZa1pHjlmYun0nSblC48160uim
faO+UMsqL/WUpby/Efz9awXcOtfVetecWS2HQNGxbAFDQlrkPnTL/OofMVt+IYXj
aDDcomeA4Tlt6qv3/VC5FSVJxezPQTCbCHwyWswLF2WB1AY47VPZk9JTss+JvoFm
zLMYxn6rFIyvB+UIESmYvJkH+DdMq1zNuJ6WqhRoVEuIhSFAKly5/yw4Xf7jHYuN
rDF2zCaPzzKISB4mHMMyK0nuik5ZO1eb17XY20KHfDiISLgYW4lfApDa8OX2kzHB
hzTovYRcQjdBssAnGF8L4W4wDbnbbbz3sPV7kf8LYpwrAyYZpVgpOuUtO9ujffCO
Q4xSStSW4qXhBdTbMmmZjLZeJZLCX7zMZiGeWYlzksaqsOoKFufE6gnPf3JUWeO4
kA+T/I+LfshWhJtJZRXYa/G5yXrsUUzUG4/JZlzqQ3iBYRCODm8FvNql35lEaUKz
vbs8HOLOyVG8KPCp5mE4W5J7kVf8EtNPmBhOGzt73M39z4K01BjM23Mnp2mKOuBo
ArBokQvGtyOIvA4UIrZZXQkKRRfMG1WsF5HFoj8evMVtVgL79hG1tfeNG1Ay6Acb
eeNkt/JBw+9ypuO7UCaMjRV0HRR/ylDklzRjJ8xkt2Rr33Eqb5Nh+KzZ/M6jMAmp
vhclGslF67at/NclfU2CkpSwo1uCnWpDRAprgc68vWO5C1pzjqFd39b8mgiPlorL
YO94KySV0sT+zG5BsbeCUSTWUeVWqV3toCZ3KWD0GYvo/q9kBALdHdN9XGn1eyfk
OfUKLcnpMaT8mgoO33wY1dd4Ynej0NmFbcchV9sWRUBTq7R6BUwNdujghI7UW/le
wQ9L0FMAr6wo+RkkgWEfxsbzTFTixt7lvh/TmoXjHDcrni3+Ae4AK4lY0E7msH3V
q35nkGVDIc8SIq/T1nb/XHLsTOXw46laUrYGJW602Z0xsVzRSMCgLAcHfDmKSD7+
ZRio+GJDSU6AB92VsJheNSysfOYROLs6B5JjzCrxuzCEMrdyXd8R3ALmOYgldT6V
v0BVSwPB2lAVjWZxrY0Q1ngHin/9wfGaBfgCM7kPr1u6YVaZxBEHmfV95sjmEPIQ
OwW9edGn96ryCHJjCNPxx9uxJFK350xNuLyHPNRhrPtL62mK05J2PDYPHi+hD0LZ
vHIl5ysyY/a9ay8UzRVvbzJD3TmYSLGAOt4l+kLxSc85bUBbN21EaMW15VfIQorI
5ieNSimoG92KLAvMwe1aWST/ZYUwpjAUlLFAhQDn87V5UBqhoiy4bINALv1RVzik
vlNRDUV2JuttjcPphsrjPO+MFL+UWXYbr7mxse1kVxsP2s8Sek7LHjeTVHJgr3/Z
JRYJ2O1AFIhozcnGYdI1Nb2LK8v0wJqhpatw1DKlMG5lNP6c9fba4aCS0j+OsQrY
rDQEu8qiy+imLJ0RgdfFEbSCs5MzvSZbzGrihJeM7cyMLg/MeLiwYbJSANrL4mMH
gB7rsYGhel+Q9KDvuGKaMzwlui20GIALoCgTXeNes5QNAmUlITwxTkQYYlQerbch
chOoL7YXgyU/YhlfczgE3ZmcaWT0aEYW2XegkGMWTLL1QUV37KFAFsC4SAP0z49B
30Pwf+TrzQIe+UmWxZLWnM6lMjV71YVJ9wJyOmSYnQZO+8VbaW7v96S6BZMYyHXh
Vv7jURnBLQ05EAxqrF722jRjYoIVdyl4HiN2yO2K9/27V1HyM4A9de+9oFhzReJz
M3E5pN9EXIo57SfnHfy5fy/O4qp92yTMKYz+Ht3bSkQwaI+9dQlXfNulw/HGs7Dd
qFAPOKSl//J8x15zDXXYoT+50GvfgJGNEuem/YaZG2JDq1kGVl2+SuKlTng6VfdH
fyZV5JlJm7ccRFljsn5afbqauLmgTAns7UIu+HrVlVbKB9Odb+wLW1wOfTG7r7Ab
6SmwkmqfAAmV+foY1NUs7xoX7rc6+Mg5AwxeoEfv/O3TaSgeboAMx5IFNo21T2NT
Hrg2Xf5IKsvMDTr7buefq4/WGj3ok+aSNvFgdBzS0NPdNRqcjcbyfOPETwxMrA0P
0qIn4YWS4E7aNb3hDyfceOUNP5lGZXVFOsvrNsSOLtHhM3yBkrZZbUXDViAt99Vn
Hj0wmoQiXkav/h0dPsCW7JjEkyhGkZAEWlqyMK5dt5ShGAYw8ysK63JP4a847DrF
ExVJ19KtRdT2ISVzWkbrIJDDDaxS8nY5dJIZhueufvRhs0Uqxsbx6q/OcDFDySEU
ggd1d3Zb+F1bzmGC1iDLM1jcVtmoIrfMqvlM0VO4JP3xN8mk07m5c5SsvfXHuh+F
1NHC3SfKjyJrDUBvYS/AHz8A6FvJxPvaIaQnjVqDAWs35hSTwTUgOtSaeG5LxtpF
go4pTWK1KWp3TJHdIbNqVW0UKTM2gd/IkGvtVVtUTy1QcLktXpO/02qgJbJ3oZz6
NDha3neGYm2/nEE0mp8Jez0zZzLyiocr6SpDZmsjGDcjfJcopGzjDRrRgzXZ+lqe
zPqaMhsn755bHY/SmLgosn0kp56jK7Hix2SwXBIvBcMVe65VtJnYBLg7qxYg2p8t
o6oeUFkPTEXYjulPApXyqeqjmqhCUT1SDm5n0/lFy45IQQ3etkVv6ZlUPkJQfx5v
gnBBNXBQ/YCR1uH0nfGl413elqnOoLtIPNodZPcsApcB6M3cL/LXvPMwF6jD7t20
hbUimqVpAY9EtYzDA331wl38cCGrCSkyjzQfWBFzZg6ShDvokJzQSN4Whslz1j6w
tn9KGHNcwzVj9v2OKGgW2DcLuY1ZHAWSiik+7Yhl7osX+MJJUv2ONaI4H+2i6BGD
AZC3Bzk/AqiGjqQo9vzS7UflzFHtIeArVqYlb9lt0oRKqnVDRS5OokmK9yryTk8I
bQ5FAVPteMIKZM9wPPlL/gB2/4hP+QcPXly7ySDxvMIRVQj4NN212kP7yLiK4WQ8
MWu/x9BYlmAwmhLFazmeqkLmZUyCU3XbaRZck7PjKufTndVDHxdWTxgwkZQqw1t5
xZZxWjGowTkj3EU1r7FtMbr/QIDeZDA1CadiG7kRqA7/3uQc1NwvtvpUzdNGzce7
wY3QF1x6DQAw7j/f6+hW2tCo8jw5Q+bY8RJza/ao0Cx1XYqTWiiGdlIgVuZcz8uc
cOqlW/zVWjQffKkj22NUEb3RBOXZ5CIVYesBNHCGuxnc/6RJsd4gI3NQS+wdD5bt
JdlZdbI5z6kiFVVaCMw5rmUOjLjmKuGvh94PGbSBCq+SmHtrMgRP+yyGHQpflEwZ
CGdpEPbYY2xtSGefYF55FWMMGlMmFRoQmda30yWMU6gSgbc6r4u6ABcLw/+QONfC
YxVgbrzQ8N6sklDCB7wwwNGC1z0vUzqAjxSvOJRZuBtBkoFXwwq+y9J7v3AY9mxl
oyV6ytRIoUNtgMaf6QSJW4S3Pu++R0kxFH6EDaXUG+ca3MwM5G4iUGnGdDYxFjTu
jKRRQHIjKk271jcV5C93Q8/HEaSu/3REUM/98XF0ogiUsStIsnqBR5N7W0B8toJa
sDW2wr6Ne+sZMsGheQiom2mIUcp7J94Zcdv3IfgnG3hqVZKq8YBHWCeppkkJ+FPU
oMMAG+R3djvs1d1ap9Qe49cjTNs9fUwvSZNNsYWp9Rf5p8VOw40LkE6QFhaT6U49
a3sjhYmtTXywN+qPqO8lDIMl2SIKXOkPz3MomaQrW5NMbIXle7TeUEdp3BYDxX+d
KX9NuVg/ZVsND76IjLrug69QM3ptR2laUD9JkaBvxwEVcijI1cvRS6S+W9jz8JvR
ajskg/NPoEOaEKnwZ1LvdbvKTVE+9r1l/acld3k73dmg+18xlXThRpUuBZUATVAX
KE52f2KfHiRCqLr5RVAPUGTTOVD8gTSBHfySis8utNw7NiI1tOAAiN//DzzO3u3t
6F0F1T3MlKCw2ZDQcQjf1ouW75/TsFEV5MBNLysgwApY0SGgkHhHBs2qSp4JCPin
TcL37j33crInkBy1NWBmJoN8nEKjV8UAAwVe2YnSmGXmRzGakXfk+ffY5Gxb82ou
Rj71NcVuoBcfprF65+B5tM0xPTJULkK2YNvi+OQW6kuKTzmEf+YxpIvypTy/HKYj
hMDt5wpuzA1GNSLC2lRFHnDwHUMc2GnQvXBjJJan0zcdyjJGo/+8dVPC4xYdfGrR
7Ekl0rkWaQOlFtNlo0ZA388qF/D9Zh1mDQ3cEBYGv6thHH5SEZl3Zup5exEBTUeY
MucmmBZp2h8V7bH4uc2YUYr3CZwtcp4uycR5GDkJFUjeA/2ientTrp6SEkRLMBtg
/mDObD4nB13vq/3HoJxzIzUvSi08Y/doG9y9AyUhAixws0TSpASFZ0/mb6t4y9rn
VjAJn88b+XDxxUw+D28z32Vbfe7dp97j8PxW+OqHvSOTB0reN1VfZg6EChN4Rdc8
1KoV/UDkZXUbsFdyaHkTb58K8N1Ci7tl36FdF8nayf16nRtyV3Xu69JxLMs7g3ID
PAJLt1AGVWDi3GoJaK6Zpw==
`pragma protect end_protected
