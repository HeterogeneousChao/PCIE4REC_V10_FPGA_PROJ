// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:26 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
noSFjPdde8joYf3rxmYH5fC3xTuzEExgPdHIR7zUyvLla0cYBz1zE8I2t1bDn0z4
DVOvc34N8tIx6sRXVU26lVgndTB5fUPhtlV7AOIZ2XcbHc3j1IXMnsOyKwNpoTZi
Fa/+8wVxu2xcnNZ0gMraQKuSzXz7XEmXDrTiEUhJVRQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
2yi467KY8ERo2BMhF5LUXNRF0Qx2BhBSvfFw+rHUQKsyVGlD+yvhWA6J7xoBQk0i
yz1iYiKfu0QyjiEuVeoeW4mFZSCmSXunWf4VfRh94Cuec6CG/UD6+23FgpXImBra
5THwdSu/OJm/XuRsMVMURJY9kzCFW6qiUdjgwdzybrs4Fek41JnwvUBEySv3Jt6s
nDI0Ixeay01MrzlseMUPm+udlO3nkS06VHWfbK9RH3ooOTh/o5Uuyo/oIhlnLW1j
Xm3pX9oj5JIFTHJZp1iN7EXqL+IUCQRMFq9AjOCw0Rt1ZKQSn8LiIn90yRJjI+e7
GdY/76P/83ut4cdS5wK52bDsleQVEToF9AZY9Zc648YqChXhsBXT3J9/rFqNAAqF
lIY6WippFQZ6qgE+meDRQcN2HYyp6aWBP1FuRcLarFsWNvF1ZhLyCqVGmvGIxxNN
nKlLtooRUT5I89CV5FR3cBlz5VE3CPSm6CZgEmVA9cgU5FGZTwrEF54gYm9EKiiW
09l4blm1dKnJjT+3w9HDaSwr0QeqOocUDEhKSeGwpCDKUsz/EM05ZifGNI4ioyNC
5bbduw5LloWuV2WotkpZ7sm1YPuX8tZ02huT4ig/2GDjesalIqt9gi8kyQbA+ezs
jkOXwgCikEkkJxjItcqGOWC5U1KsV7Y5RteybF2kpNnd5Ht9MtzfTVtHky5raNtr
p/vJWy1qh/Lia1ePryNNx1y1W4YAdgy8pLiVu8ePd4XkFqYzVc4BoNOW3uor3FHS
l/qsapjTzvZGDOwd7GwlEarHEsudwRi8Ttby5wRbsRbtzS88kdPLAAeHnpg4kD/P
S+JGsfnOwvtBmiaT+LcbD8+brLcV33kS3maw3nSxGMBuwRP/bd4yAMYyr9l9meBi
HHlouUF/g5zRRsGXddTaIzjNHWVvvnAdl6nW3Qrs7KP8oytWvit1MwNoIBHAhHWx
eiJQ6YUdJPMjM3MgAcQvBjB0pMrcRoUrPd1EiGD+nlef3R+g/E1Ez56l1YTLu3qs
5LTmJfVwSvhFPx+HmrW3CaIwzVA7BGximHwN7mTnn2IPLYXVvxwWoKxznJQD/xsK
RtrDs8+DFHmy1dDhYrHeLLxLAyPtUfjX5768Hv3JQfjZvReasGcZir457IpV87tm
Kk8dVgaHGR8c2QcvGzEa4AMKA66Fvt9i4SxYtFYbkpq8IkvboVW1u67Pp0pmORAM
BZmmW0kfkFQyb/OTojK1Xfhjxfa9x5ENqpPliTMAexekJU/x8MHeeB0tEWMbVHCc
4QhDePFh+uGrKRapSJSZTgofI2F7pwi56O/XLqeLSPD543fVd6GZjJDVJuyDx37X
9h+XWPG4MN0xKhrn4OeSaOizO9Wm7eZMbUIetJwlcTHvtwb7tyhx45TYTAeIhZpP
onkkSYo3v1DS1s/30/RyjHNqPq/ghauJuAKhgogyb/7SDNDxx3g9nO9tDE4IO2r7
dWi+Jj3Y7pmIoWyS+64qRD3y6odQr3IgB04W+wzkOjbMsTscikXZ6QJT68xalbHS
1e0+N+zYDp01zI4zp98PqaaRHy9DqNe9ITTyGNJG6ECz/IqFIkNmOBBFWpkzK7j/
FhkR8arWh5hWL/5E25ZVXu8hr9gUpZcoG44wyV3LVtuynwTgDI07Sl4BTYwH791q
QsFBv/aeBWOgt9aJtUOXdjBo62R6oQ7a9/s6xkxjYvgA73Eo8Qqd/MFGXvZ4aIw8
wVjxVMi85gACpNQwEbW87KQW04nJfxbcPJaLIzL2Bi7NWVPOLwsEjmfmDd9xEKVs
2p/uLduR0nB6gTYVxAmOyKmQgKVISXsyFPOwebuyj8Iq0vEzYEgh7fU8iwxanEQP
Hx5fHN6FNtmFGQ6vkTrFke/MXhdzDwOVPPQ1w5OMxe8fHZ/xIMrgmqfHE+jUGCtU
EwdVGG27x56VzjLihxYOX5BzzQiESZNDMkpDra04c5l7GbnbAXc+Ch3wvPTS1UgT
g648VqNHrY9KZAYOoGrSAyrbbvAnRlvPGz/H37r/t2feNntb1S9Z00WLl1x70lMQ
a8+GCK36ezYkd/ozAm3bM2L+3hrbxy+iwrSdDkkUSjQdVq/sMXqC5TiRZResef1A
hsdj8qFipFHI47yozkBm37+rXtc5iv+EqExAjQF5idaOe46+BqMKh61mcZPMunKU
1xgo+SzJ3AsRDk2dPT7cjyQDKEPkZ+wxTXMdM80HKLVU5XyLEVMw3KDethkWg1G6
2Kf1NkZlZ6bZfwC8yEGHDAM0PVZh8+fCxP7cD/Hev0EEXi/lbxQgwgzSoB18nUF9
Fo36cwaX733xTdZhh3JiTOXd1deGQHhBIHXE9sDidMewq+GsAsS3stVdqVfd7CsF
JXSlA75AJ8b1lIfANhDzJaaO2cKWRmavQCKG3018C3NolgD2+VrwWvYiiP7M+VLn
j68Voih6lugYnXDtVYqn2cj072zDKHosoJpARx64zH2fBb4yYszjQlq2kDssFGrT
tKskviNk2HyIM7df0V6PrEhgceox/rXC0gskHtYwmaPYQlyITO5m7zSOpVmBX4TF
hCmuoitHG+CB/HUj92THKHEax9i7L+zoiTHA7G43NzpMfkIcnE/QK4MFhAlf/yG3
5ACgOglKvD3RJJUEFtiy2IJBP3WNOP1Qu3juycm+oJAbrCrjuUl2bgRSSVEM2geA
6COE5Bc/2oKrLdq9kQCfjtj052pNLxGRE8f2qz0xVpkvp0RtDnR23PoZ77KUcIP5
LUXJGkqGoww0emTVADWOoztDTQ27ebcJN2vm1KibIw7aqWgwC/dvgPKfp/bwUbsh
YTC3seNqjqeDrRGdYyyLOfqNfP3m5Q/7xw+NXbnCO5wY19bKQ9u/IahQm8OnbKEV
+rO38wGp4hKFJpQjb57a6AfQTIVG5+pHIru4b2hYklDDR7Eckc0NTBWQ2/yJNqGE
0GSN5hLo79Tx4Ecub4wiP8t9dUxuOxOOEDjGqmpMNUCS4ehMwDm/tDQNFLKWgzoh
NB0YjRKWiBXfjYIFksSaICuv0tuuOAm2nKzoDkoi5NnqYjoTA7/AliOZHZmgw6Yu
c2Ha7d4jX8KxcQAB0GZmxyl6q09rDB8RzAfD6xER+7A8phSO1tJL5chacl6u72Jt
3dILOXbcKE3xTsND9S7FEPBZMZuox9o/c8akOSjGXccZM3WtL5ZxVvcEZ8CSjiPd
KsNeqFTRc95lih/us+De4Bdq3abFgi9M17cHTiivahylvjbyZ6k60eXeCMzouGBL
5mfaKWxlS8pUvyyMyJa4r5ACWzr5xb52lDq+Si4eW30WQSU4hHgvPIs53krCieFy
PJI1D79fQvLRt4JVwJskpNYpj4edQzUGJUitWPbN7fo6CoO0ZfIQBqiX9yGGF9wy
+ozgZTor5ODie8wIcT8rtDDPv9YcXEuNpBoJeux5DCZllGAs/kcVKlAhSrX9kiAv
AH094ItWa+UViFcilwAqsbMrQyFeXzNPv2XkE5bYS8lRVnEnNMqlgyT4awiu8S33
soVUda3hQ2DUFB1wc5RMPefutI149r2jjosE9tgMjEK4XB537wNHGBAgeKIBpXnt
DE6SGxodnYb0PuUIog/LLRyeDf+TQ8qEb6cpOazlC56g8hmsFwL4wNFe9r1wJ/Wn
Hm43xVloH5njG3dc5AxyxF+dw1KX8qQYPxWXqeqGJtHpsd+INE8slHtDGc+tHRFj
FJ2kPgaVtAS76WU0GxTKUNbKyfEZN9e21c1cmDci/3eT/NV0aNYQtO1Q77PIHUpV
jjDGlCC5RKT5MGdoUkq1PTOZPSXHmM3e+928DdpwHTmXrs90bH6hNlHOMk54+F4t
tmTXOcpGTTqeEkkz5/ZEK584+aWncb3tOcTshofdNXzPPNrnKH9L7XXgvCFRRYaM
ueTJ+wvk9VPVKWCowj0EVKpUNT4ksh6mQbeHDBm3cCQTBuu6NEdOtE1opsPOLU7I
duT4g/ryTvTjHz5/jfIRFqNoWFhW1W7krWo1by8Yd+gSsoVmAWm/FJx6jii9xo/3
d+kzL2pQubf01ajdZa7H9l+1I57H/gC2UnSvY+wP8RnSvroRKrXPpwk8w7CSPa2L
p3TzashpMFYIYngdtTOd4iUzJz48/HwXOgj9ZiZzhWovFdUfCISCjWah11i/QjVN
MgGdE8fbQ2t2VYowje5O8fXXBZB0qjjR7UxFxI+hxvZkkJ9XzbmsIgCrdlF+hFF5
+d50JL0uTsLIrgo3vHelmRhFfG0JPwgVGSBudwLKJFKjkoO2HalrOyscWZgevyHZ
NvTlu8fk0lY6YNm+MoexlfIcHfgup8B7uOIbCJ2w3ldOZScTWZ9X2OfCi43LKpSN
/5zcO7DVbRY6lEFgz/r2OpXk4k0CB33RFk3tm9U/9JQBJEKcoTgS/xHM9NLlal2l
vuHkAJyo7LMl6AnmLD4K6n/4gItYVVnjg8qOfAF31AP1WQfhcaOKiEZvEN5vV1ff
wzg4U+mQEgLqXWn77phM/WznPPuAQ906sXpfc7fUw8xk1CeT8OAmuo3OBFyK1xz1
DRAkaWuevUnJ2oNsMEC4cufbzVsZN9ZYKFYntSdSDFv7nVIB6VOSqd9Fhe+V0G4o
4l4mCHwAOUJFNhS1Yr1dYGDD5SdUVuW3OFeiQvvlTN+/Ug8iQmJRwlGZ06OivszR
aSYc/6Td/kJr8/nkmTokuown8Fs87+Enpal2xGS7R8LpXlJvz8zUGEciCkopAeAr
nlQkaRWy1++pzP3sdQxOUMMUAaKz5+dS9kH3oFFscsO9D0UEPC99Itd5IKAOXu89
TxvYcLs2UINSutx/YmbJs7PViMqQI2iHlpiQyVPnjgSCCaicLg/NRG4jfIqvn64q
RRty67+EPGJT6lUKHnHsew4HReEmUIpctB75kaKnE0lLrHjQIQgS9kYhNJlp9uhl
ok6AAEPRqWSuksPJcYipANeRJ0Rk705SanE6kUazbQiPVuIpEOxw8CFST2Mh1xQO
OrWsuP+Hk9DxG21FsSZCF4Nol2f9XdeZUqBuqcvt6npGLtJBlbKWwf5yI3p1pMAq
A4FgtHjBfj5TFcDIXmP/nsJLT5r84oqHz14A9OXg/nsEdTWOgr4g2VxcrP/wDiNm
jPIP0ELw8mbsqj6WiAlhrP4VrZdzT1HxAwMqvJqXPZ/XXUEvRLA8/28z7IBhEEuj
C9ra2/tuRo5A43po3uA/Fpe3LLlGSZid3EWj5AlOyTyYGj1Cqmoa69kOY0Annzv1
Gvyc1WLguBe74EomO1F/EGWrxR/85ckQ4PFANGoBW4AtJWXyVF0eSnu/Ebe5I8VX
bXuQUC/qiMQPXWQCAXNnW+ioO8gdQu9UJsNshKLCdCoi3UZJpJUSQUKqfEcXw5jM
acS+fNsZcdvX4D4fEJWGDh9Rezu6zl2Zyskcvqqq7i78NtvHU0IZpO+ud0BoGwLf
TT6X1m7FXpXf7gvMdY+BcXC7oL4jVhQAztbetsh6cg9fh3dQ+7t4ESNy446qdjGL
ptXANwIF9wE4mCJUosqcf6i6aY4Z3ZJzIySd/rBmebOEe+RCy63VenLM7RMb71CB
S7+vo2rcNw64QmAouslhfHViTeF2+FFCCEWQN64bFgIa3Pty3z0gafEFKl3FGvGC
Lyl6FT3aiYo/RQcYY6QSmZlG8rPAPZb249xNF/wfwLcjh01+ZZNgYtddytqRVxvZ
bvQc6ev0/w/MuR5hwhDc5aQgoQ7kX+Agxd3Oyc58/N+7REbbVmKB3O2+XDnjZZNK
V2pzkPUCZ8G/22AqDeUYfTtNK+T4ilGFaWuYOB5k31FSfRJF09TBR5bPT8jI+wFA
3Pp9pWAL/g6szrabfobvQ1sHHm8du8vjBvFUAh/rq7lzWWc0yVXxdZqnNFdWEXJ3
M/w4jZEaKQzrIsYl01XnmDy00QekjkPLULrMb0ciRGjr0y0nldiuFh0uKyh74ogl
PwpxFMgSYf8e4WRIPjGH8+02Y78PGsWar9iLlqIU92STMExYMWuhjqU3l6WP06Yl
M3/oqkR0+k2I+XEF4FFJ/WxiXw8jZweVNaYcvKfQ6gu83eHDY2l4fGs3IArEWvvP
Gj+T0Tdo1VVJ/9v7YNV1+XMPyAkxYUzQzrT50BLDGfCro0fIYyrNb0u64X0gKTdb
kLOte24+hEFe0Si5wM05qcDPrNUG1v0kVvGx+xtFYa8lzC9l2pHGh3lEfvgS0Tp8
8IjB1eV11ymexljKT/pId/aTyN1z35RRdfTfGeqWUJJ7/GRpb1Zd/GXPo7Y7SywQ
wkNb5c0iS5LP+deJ9PQsJ6u5nPONZbvfy6Y+mE85vHGw7aBY4017xcTSZ22Y73cU
oHMxcM9ssDaL4XDRFDjhfaHXzae+K6yMu6RNDdlKkf1DstrO5SAIRcYBODlCQ3HL
AfQrrfQVtR26mhLVwHXFwM3b+zMDMIUOoCXGlRmQniyDWAX4F2Ub8N2K/NyP89Jb
baTQk4gcOLTnibFYoxbNrGcesJm7bwlhQvo1n7QuFsWOB3MneXrWZq2Q/j9f5cw2
JF2MxDdEhwzmnbJGiElAfv3GTpsR0e3WX8vVYEq4idAH1YKLjTu5kFtOMF0y5nNm
aSLNcc1r3IXc3EMLMf/PUpGu96bHzrw1E679aTH+QGLT1S0vwdn02LLhF2OaylMP
QpxdpWpiyp62FtxzG9FRg+BB6fUW2NJR1HtE/AHxBaNtcAY3uWWJgNRMPHbbS3J4
yIcslAxv1/q6nAizHndMDsvRGr7SN39U5ydCzIy8hLBdKtizOWJm5T0jb92WqD9J
lCanJJvZJitWZHaFu2zyHS+jGApMCYqaYV7UKBVHd2paVFgA4ujy8cRv8456m+o4
abr9lgAwLFT0GXbHb0mX1BPW5CfhWPC4/XyGvQY105WjjP02Yn/eR+lvKPCj06ct
FQ0VB/DLdph9jfHst8VsyRqemMccDWWcT+Kd/8XA+1vtTEkmkmzIqVRoi8JLqXsg
asm4r3p5yf+EcRDikJYurHr5MBJ6LlgaMTY3xFTER6UxvZc2j5cwxVi2mG0VSKfE
zzEr6FF8Mimlc/Jg7mdmkIALEr34D8DfMdR5uipjhZvwpdkeIKH1KIFqV2T0Jx+i
EwZ7BgDJENYlUbWITDjwsiKq/jU2HfmHo1BCSPYeFl3/W+bmiNA36Ndq7zwz8H77
1OAvrsNi9hzeRX/TiaIcC3knsS9BmJdPOmBQLCBToHlt/ZXowiQRdOcnpNsqa8MR
3bRynsgFKqDydEw+t/NyZbU4FiOTg9TXkqoMFg58HtV6Qxw+r14mlW0X5fPEjKRh
G4W6BoXxZzIxjKW+ztp9hiZ0bcMKE7CsvIEXHQwxcIrMZS71kwa8r593XIsG8fJB
m+vpcFrFEsMEq4x0N1dBG3DjpbfJKNAVMGrsnLvnnW8kYti/Vf946EGoRHv3TN4V
rrnj3lpvTaGvBpdHA0M4wHLozSOCafGD8Rd1bJ6mDjdC8cHMZJSapZ67Sld1ebhU
iFj/MoLXa4dDsYtbxcumNNQKq8BkyuW6d5cZleb/EuP6/cy6k/h7D0lJ6G4h+Ao6
PATO3w2xwoTl2qsU0Eni8x37FAhs+GYz+IBnWCrVAoHXLDq0kt5vqjbB8ZKQFvBl
wajXaNLwrOGakCtr2qVLUJLWyEgxkX6Tuyy7BcnL1AcswVvmj7Gh8ZgAQ0fcixsw
WDMEyVtWvctddFWDHSfwhkQHUWZR/kfyv7KlI0EDJhZlY6W/2SPk3cuN7/tWiIut
vUJHSjM+cHKIeXp5JURZUIZmL2QGLs9kRQAVlzxqarMcd66JpC3kFDjpFFyjLxpy
4AgBOkcJ2Wf8GyAH0x6c4+dd4dDmjS3GSGTxh+BLzzcDbtglO8u6w8BzOyYtcInA
Ma5ScJLulCIHHSw6YtNWCEAqO6Hz9y+MPweyxj7E/LTEzoh0D+7TKHLJ1E7DoWRO
miGCtBoTzBgqT7plQMfZad3RytuM9WR2pFuXWEg/sXs9Psc0FDbapl5QsgGAcvF9
yTW4abwMgdwp2St+jEhNGCC1vcmbSpht5R2E1tup2DxIAR/8VYR3Kob4jbez3qHk
EgJlqFYtq5mLrTEiLw2TqKQ84iH3ErdMmka+/WEq4wVkJoQqrITiPhLGZGEz0MXQ
8jAElchHDdg6g54yP1kVJ9KkmPSDCHv8T1rhes072L/mzKJYeJMpEaQP0pZ4MmZW
nvst4kStgJIwKlQ7+u53dFeKWaaevJe8g0Q3fU4eQ5DBMck8bCtYxMZ638OgSiGM
5pKj5R1Dqk1rd8z0d/J2ydoeOOtttksE/5n9JVFOAXCKf95GVrxKJHYWDhTo0sEC
7f+/Jc8uJH+vx8zof2PT6orUDHxuIwKO3s/++3pYJITj8ha8W/JaUPWwSh0BDD2N
lv8HDDSapKd3ZNtsMHPqA5QUeOoF02dy5dkMZV5MD8gEEZ7MklUEPuxEW278xPr+
Mbdb/4MZmdNFBjEbGzxf5db4w4s/1rObBIdYUjhJ6uz9RUyBzxLZRdbw9jWFXGEM
CizhKNDvhgnWhBnbIjMzUzf9f4UX/IHJeTq0GTYgrrPaClzqrtnRkgZWWi2Y92C6
RaGaNCNTrNPzMOb6v4WhNAtndHYK3MNfX40aiJS9cKb2KdGqliyagb+9GozvbbIa
3sOSZE3FVwp3gwNfaELiRRnO+ruJtA1ZA4+iIrYf5i5hmu77swHnFaTRJU6z2phT
6sOutZbkbszX9StK7ucZWlFYPY+3Nwvlt8Wvam26FHf99qXWLOW/ZYFqO9hYghj0
bpIE+cbreTX2FWQOmCxTBpGXz30ITgjF9xEj+rWvnix/sp0uwFN0usWJhBKXKPqX
qU5N5nnefoPWue5ANcHz5nxxJrgr1RegaZl2+55M+dTQRYMSu3rP6B2B/Y7mWeNO
DjanCVryfAnPbnYgAJJTINL/ioHGy/ZK74zbLWe/Ig7TF9sk+ZXem5/kdTZdDCKJ
hZpwFI0C7EavVEEUHtsbSoJNZBMY6jStnZ5zlftYwbZr0XZByjNlc3tkfO8KBUcN
r5s6QDYhSXJwP8YgUl6Lu1Djv0wN/SU/+xNYac2StvWyyyHam7bupEGU7rU80tb0
SYMJ2atbADNlhI94H5cO/QPoBssnQsQ/8Wev1TCDa4WbzP5cmO4p8hBBMv4fMKTk
e6IPxdr/quMKG1c5ynul6Ep2CGLe7kQrFIAtb4dvU3cHrKC04GWTkKYq/Ukl0In+
t7u2kgXjHuMIaZabS608zC2JJ4DDwqklsP+WUv1Inh+TcEXjGuRMSavehL3vnDPu
qRrj9FploUBt4SJH0zFj9dPC9AlcaTWIopz57fF6l4LvMhfEdY3qCUvIJbYS8MqD
TmVfo60s7ligz5aFVrek0moM9o5VGjTHlsUBMyh2ZCkoxAOwPOplel51gCiwxFL9
+nIwQ3y9XYJUqTPfsGC5WCNT/PvjNGFf4+gMUwCLFZ34UpgfKwvyy3F8J5iac+Op
Id7Z4WVsfjccP3HxrrwDmazRMH6/fDnlqok4/8ZKkwAxFbHcPxDAFWUyx1Tfr9oj
9xMsiTEiRvzo9on93Yz44ACPy5cVZVjKOA6A2lvu7FNBJdpknAq1MJk6oZVd98VX
3sH1FnGuk3pED5HdrJkKARsxuY5H4DvmrLTa4fQ2EkxyGOh4ycErM+mfjrQiUn6F
YevrwdMiC81UeECvBikKlWpwfX3yaRNVrX7uk1SvZJdBw86mSDM8XDmb2gza5t6w
+w0lQBisAQVlDruo7W9sIs2AESQm6BnBRyBcvgQltmRQ4tZ6vZ4+7171NWVGTEX9
bh+K7mMLUcQg/jhBHv3+RXLGpULk3Yav9aa/BznLZiVDaD+U1i7zEHVepoYZE05E
INxTlZd+z9kJ9dwv8KwT6lF4tESGaDFK0/S/IWcZK5y7NbSAz6B6QYvrMNc8cnJb
FFkliMM5EfB+OhAV0COgH7KRfv6AozUUmCaCvhsQg+fEycTaRtrOdV6PGlbBN/E3
CrOyXLeTRHuMSB8XxZSGjHgnLPwyaUX9lRMWMiHfM6E1eUkWl8u+9KXsYf78R9I4
5MsEIA/Io2Qfd9n+h7kOoYlh0D5V0EDMltoMNp1ERsx5mtNqXQiJuUVLg4vfwkdq
lolYixcS72IHDFwylGsHVpGEc5H7cwyMca+R3CNgJ/V5tUAkWJkpldS2D4F8uVkV
k0B/IS4ltKzHEnhjEZ7XPTEI8InPsrbD02kMp/PYl9DCKw8LzU6gjEmlL9uD6uA7
Xs2GGAfkkjVyTQtIgA7VUAoDlLlL4f9zjlO881BOuP4A8I1xKFEOCf32C+e3TgS0
H2dM0KcqGaAjDRxMqACSTwId3d+4f3irtAjBEs4U8MOJYyAZDDuURtYTkO2PUuO4
mwFXnSoN/XiZVxbafMwR3Bz08AOWCMR5+Y/VlYISRxZFN00c2aU2EHEAA7i6xnb/
cFJtejzL4zN9fcEbHCkXC9qMTSp1EMaZvjMQs5yKsVCM0nbLtseDbeMg7UtB1iji
N8VgiQAjJScZTEWQuaKFC/FK/rqy9Dbzck/uQwlK1VqCkuaenUjSuhfAGlCbVNOj
+gXqUpkbO9woVOtvY+rOf7+agCaabHg3SUYyw6KrxMYRBrkFIo3lVWAsvio/A4iR
lVQAywQH6iVgiWiZBLLiKg3j7kY6tk8u17Ajx3RMIH4Xv1lcYm3nDzM7eBM1//gj
3fljLXiUUsmQT0t/RPEZGuGwWKEaqR2axS8Wn3VmeX/kP/VXCYstcAoZDM0vXDF2
J7I37HnIr3XvZkPqQ2ERLAFsmIUvaNfuO3vBFGAR32W+VzFpwIHtMPic+TiDDRIh
gHaEIZ0IJs1OYk7ag0F7lX/1QEfAlMJyobXWm6Jklre6TNwYlXIStYvITa3if4ec
5p1Z0+yVuiVgs8rgkCXis+epsChdwBGuNLqksCrlReqCCGK0b65Zgwh4yrTQ5tJM
PetVSKAkSRKAsfOZBN+iQrx1xn9L8pC+wsVDAZkpTRkROWQDMDdki/gCjdX3OViZ
udWbGlpP0IS9DsuIYaqBLCJjsU7r9cHAdfBbjVlKGhuaD4P/SrT/2d/5oKZcI3EZ
m9lru0extbpM0nofkWLjZ5jwqnwjOKiqMOECOjOs+/sx4E0+LQMXDjLXboV+gsvc
3bOwgonkHBLHfAgDAPtzGigDa4RY/m6kuvPKP0nymFD+AKJT2/VJ4ZSfJCDJBHGt
rKZhXiw7waRK3/rl3wVjdTdp/i6+1RnWwvts/IwUT75Ii4r8BNeLBEtsgboKCZCz
WPgeLxKd4Wk0D99LkNahFUn4zViuQDm5a5RgJGNigSmBliLF6B2++sC5UUd6he31
TcKfqm99L3AECAYChaRW6LHC5gzkAC5L68WO1oD7BewvTpUbyqfAWb3aN6CL/fHM
jFDC+1UYUmZGWl2HYyfzsCfntV39/KkGRJKNvuOzr9esPm7LpQXg+jpdXyI/Tmi6
eBuFx47NOGw6xi5hOeDX44n8Lcznm2N6I5EmNoP6+ApQ9Af13JI8GGbWeElhx492
HJR/Cr9FUr5rAxloKGAD3StVmwYNNbJ4tVBwQGtlYn/dyqZrtepT5gmQQKNUo1I0
rCWrVOSS6b+/hs5GEvtxFiXE6am4hUg2HExhADbyUwClCAeRiYlGshraqAucCigN
VFLPiJxxHj37JssgP6+KIKVBP0BZ0ie4H2BsZScv9RG51NQh/cqogbRmnPIz/uRN
Q/SQNfWPR7zDhaMvCf9+85WveKFFnvGUk373w7Kgeuf2q5YEkRwmvRfCntDeSPvE
oqMoqOziSoDkuffa0KVLtKFUQ6M9GipUqOsLb76SUUzAq0qUGV9Bm4IHtjb0l5lB
HPlCaBmaya36X05YuYNQiJnL6C3fwkNemDrnybzNa/7CeLXnB3T/QbcE2xuMoiAM
Rw/Xv62OGPZ0VU6zPbgHhnA9iJWpxHmXwaYTL0ljVJZZNjL8B+tMDhiaXvTZN3O3
KKMyf0Jcym8drV9+EbGVYRPvJqaC/7IEWtt5k92LAi8n8s0bbnkYQwBFfL9liyR5
0ae3W8l0JKlLP6Q7lrnOA/gXBXexhBSBzhCloDB4FLjhF5cy3x7+Z2hxocgyV7z7
qg7G0zITB+hoiJx08plynOXFpINiV8dt3s9meShM/9u6HvpippnOsYeRFyhB2bQk
jzk32zKabWfzviHgBsgp+vXcUf7VI7R1LPZhgZjl99IBiiZL3B8ep/7XwCfuCp7/
WEjZVYe2VI96CBTmlkPSrkgk0koOCPjzeqK+RJoTBWFHi8xECXvJB3kGEWaJGfB7
q34+YgOrVBbykuZ6OIWuKhH4zFMctSVexisErZ2hAEAeKxZ88pvp4Sh37KAujuos
2VsCIUYwXMogU0U5Hky3MTwVf5qMGpWn1qmTw2M4MhoMtNQrIrZ182b20s3RMpAt
x/W/gykzCM8WqaREasbPbZAoE6DbFOMnqWrQMcg2suYpIS3BtysqVks7Jt79K45m
WNdznFd6AE1kMs67UJruTx+RLKqGNAyHj0D781ExCDj8Yr1mOs6oD164wFd5iNJP
pcWSamFBimlKbgfN83Cdp+dqw6rHaaLYOnTZv0IOEZR3cQMBhtMnRB7ENV5bmu4k
ipleTRYrPf7L23CCTCvgk4ChCPsYV6JUZm4332TdnmXxE55uSTYb1gIOyrUPKxa7
C05NKO1qBFX1EP6faizjtR/rNE7MVHjfv34YL+em/IrWWBqhGjYVFfC3Y6FThmri
BGxdegwLWQkXBK4E07/HY1l1PU+tNNIeaUgdeuxQlZtXccDgQYLvuq8IM5pqUrcr
jTiPpGmVdeYiLSv/MwOAkF445YzsHHBoH+fybXtZqvmZDSI8b3WStNMFb/8TQos9
Bo13ABwdsZwajxmUqgeAyi/BMHkmv+ODn5wB0ykbvz+7+/UAT+RaF0WlkqE+0Nz5
KHKvVORGpwpHcFrZkgoSIVio1q70fIK9K+HTk2EdvwKTugtQIllVY/wCJSxW5Svw
EB85lb8AUY0VvjypA7jfPU+thcRZSdJDNup8QBKkCam6KghqP70MdwwL0n7S6ZEU
c5KnCEOIgdNB6YxxofcB/85Hz/atts9wjddSqdog8aU8XMk0cEFbIWmUFMHbeR4y
BmYWNnkZK0hF1m34vu5DcopvWY7opPdNC7phqh7nRFy5mnvJIzGA0Jr3TWBsPRC1
cDxTeJ9hTw+LadwU89jFiTmRvEum1oHaUFfnrHGdW1ZlUhdF0T5Ur2U68uSrM4pp
sTU3CsuY34IbT+G238V6D167s6C+7Fjcm/T0vpiPODJtws1zjBloqZjybPCGIZ7u
ovqkJqLMdhCfxpx3q/pfnpsKc+Fjihk6PvchIYRRgSNa1dTMNEoifAbcQc3Q6aCv
Zoy4Kvnb0iQWMhudXTOSfaOeMlnKjSPHc8jQeuzkqfJlymUwz+v1i80RYXyU0sx8
Tq9s7rvdPw6th32dkOOzvT7D7rHsI9pJsWtHr2S0y82B+vpbeItmk3HqnipxhMqp
oOmOsX+P7ZBoGjkvUOXSamtXo/u7DvknplPTCQSkj9UWgpOCQPD8y2nH7YAGCwGS
la6oYRLxTuJlzHyUgmVzp6q3OILhNzOF7LWMgn8bghAzI5uTO5wL66Xuwqocb6H4
HAL/YFgL5IReLTB7qunzPDvkl3+YHaBixOg9ww2AOjDQjWYC1OyfzUeKiZ/CAMRV
Th0nr3v2h0NYXPTuCHrJM4ZTMlUlhRuSBFGSTYqgU/reXTz2XMRPk+aM6xO49JSH
zg+/58nq3oIbovRaqmWo5N7youRCwMmar9HVTWx+37+HQIl5Tmhd2rYhPXpN+sVj
ic/Rn2BOBUj+RIjsLfi78M6RNC35cpgoh3fDNi3TzE/HzaYPdou7if/EHwRw7e3M
fJlecAsVpW90CUZb+TNtoel/i1Fcfirqs7gJdDSIkvlRYPlf48RFPYHFU+B0Emqe
A+sGlIja3fJ6fcD8r/f4f+OCNRZ45fZ3alAKaG8CRzrdnsB8KBmSsg6eWPT3Klwp
ZkhxROgxvAr7uX+w7SuBweOUOLWDPcC7ZsmdurQ+HQugixbGudgF8arWU3DZfz/2
vAv6g8yeyL9oYaxdQOZ2gV8AXWMiaVgS8/MhVW+OUbaJS8XuBK/tK4guzd+LkVks
2t/USISAvKIl7sLvUCMAKxbkAzHAK0zP1KsF4/KABsiK5H/eoVR4I+hdSj3dIVjj
4bTgETFyaOgGl7sgiWbdBeGMSIkW3caiVrkWjLRy9ZrGIUFhJjuJjWS0IamwDaUc
ULc1r48S/5lEQmtDeFhhMpYy22TIuMdqMFPU5eDFKrhufDWdXWd7xXqj1JXO0DXY
SQoZvXnPXsQ6+o/lH3HKXgKC/PI0flIj+sWsv638yYxS99Y4d9ok2r0F3A4/rPCS
cXLwLTpvVa6vlUqkz46TiOZ4qW1xH0AHoaswYUmOiGZq8E5e4HjtEdKcLFRe4zE/
4cgblmCjadOxu2QzhG6GP73bYddBIzuYdIFXfFSCqPwwXfC9jDPv+msOBrCCCvmb
sAVwsFZsy13luJXNSED0FlzOXKI2bizoxYRBsBLurIeNxq8OX2XVsDxc5WSPUF+/
BBW0kzZ1m/BqVmW0dOg3U4D5APNWGdjEaMr1dab6AjRxjm6caTGS4MZHOQP82uaH
ijPsDF5O+otVpNuTHbXrJISbaS3wn93iWLYF082ElMiIcr+e0HznJmPqZuaE64xk
ntykMROWsr4wnV5osTKILu2r8hGaSzSgLZolhfQLSHfb0IBErRAG36jrsuhmgDwE
WlFxd0z4gzJPh/Ij9KtwZy7PagSER2MBpL5zDpeV1hUvN7+HK/1thZRDn3TxL10+
tQMoMj5rUkJ4OtkHZynspoeZEI2Ivl22M5SzL8Hotlmxia8XgxDLFmdUgomuHh4o
yGttkyWLAJFv36Jrgz8c+kvz28hfSJi9O3ZucPhOyR6k0infpbLvkSflbNvDaRJP
5Q8pAGLKTJWQe604fdhn5ePH5R2hYB1GomzQ9WBKN/Pdo4XtUGAk7KHFMYIjcFoq
/on6JpSKZBt0eCV0MzhHKsHdPe3xj89dD6rajc1FfoK1yCCHuz5s2tjouEw+CTjS
0o/REMp6d4zNALU/zAuFmYUwWdrDVm0yYbDQkHWU/CkAK7NBKXrHwC4Hbjx8UWO+
fo6lc+g7M/XmG6fnrB4IlSydv0lpRgsLbojL5BYvYSepaBiTCssdTggaTrRbaCpg
w1YIconElZTetQBt2Upu0UgEdzMnSuokemcozwh3N0qOFrQtDfCu2dO8TFwW8803
gG7l3KAgR6+bpc4Reg0aaQ==
`pragma protect end_protected
