// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:27 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s4A3th/6qiCCj5oSNfklXXkhjQOv83MBJ4m5Iiz0mR0OMUgBDOglZ15nXQmbmIPu
+LL97qC0A2Ypv3pJ51zHuGkS1WoGOO8Bk2O7G2jKYCMOB6fZPUnE1e+9DXC7tGFV
QTHk0UXt2ubekRHr/il2FMESzxn9bqms+i1mANRQHhM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32800)
ek0+f4zxALgyO63q4zNmxfG3/fQy43cjDcJVGi+0RYCTTOs1AXnQIO0UpSHpmMBR
svbBK25WpghiSi9WL0baQY5CS4QpsxZPwuFyJYLwtxotY3iABBv9I84+bjWCnp/Y
HvFcLdvIL51HtZNiXi0HdaIKykunTl3bF48GMz6Y2BB95qFxqd+8OGVnKLec8eYN
+EA70BlDeACSugpxgFMb23+tDUBdAk6U/JHvRjyW0rI86X4RaruG9bNmudrO0I76
utKnO0TXV5/FNqTQpTP41TQG1wqlVcJ6bMvzOkqH1JIDHGgBuWa/zBEc5bvuv+uu
BAnGn7kdxrAtzT/rqZiLGsrguHDHsn5bEJw5lJuGGM8le+NHajLnpWUF3+vl67UW
0wfEQ3zvKumG6Q192QDF57mfchCyI5Ky5P4t459ju8lmBTIjs3ZrVwoPFuXlAUUt
1KOUu+GNt38MCj80Pv8lvdFw1gNHOs23E5p7KXXqh3EM5wdbU7UAgDMXC+azNxI7
JsmzHt4SQa38vpBOh5wcNgL2vF8NLvi0ZUGlRM+fSdRLfv4zud9CgVA3W/bmvhP2
7Y3qgWpdWb9CSFGWZgZ5/WWjebI3+eDYVGoLKdapf4EBRHpamQUmxK+gvjzLRhcH
lMIvJnHn2XB0IRh+EIF/6inR/l9ub6L/pvRX4RzxBa/0N8S+IdfyxKY4GR8u53xn
ywfULnjAkztJKAjEPtkwhRB7d55rFHB6eSI3OrcDLnFS856OR0Tp5o1jCv1q8YlQ
YA+hGnab+Ey/6Y46DykIiuuymOzN+sH7WwsUdg6A0nO+DQ/pXQWGtvf1C/hBQspy
VNovFDand3+k49vBOJ+CLX7fwtXUYfHPbxaXl8yBJKhtzBpfH05lTLV4328IKB0k
OPJrVVVzaseTMjTh3z0xqyT//a3+Tp+u7tsLLY27s6J4FRgv9NFWk+1O+4o8ATZr
/Wr54T7tXgwUJyLa6rsSItPpFMO7QLh+hykWhdXFRFHNw1XsT2TJEQwKE4lnjsYD
Y+BLbArZz9eQcbVANrFlcYzGqRj2bDqIMI22dSugaIcs5xyhhGk3JgmM21165Vv1
TG7sWcj9LMghQirjSdUBFYI8t75p9t1oOF5MKYjcAnK1hEIGEVqz71Y3VimxqF/j
PTNt9CdKU3lZu7n4v3DM9Ed3qJd7R5FyIQJB3BHPsBWuheUi8aIWNP+ggBo+sTPx
ntWmdToz5gp2IB31+XAdH/n3HrmDkLP+knxE/UFzr828HXQxfwRCTunBvttN+NQ4
SgQxSFtaCUo+VHBdM2jfw9E/onWTF5TVZWDzxSgIvMvL6lgzqMjdMFNs3NbHqzS3
0XVsYznFex7M8x3WS8Vx7gRWNcU14fY3KHmAENqUCe/2xyZXFXhT4iMpexJSxbE7
a0bWqYn3bYMAxZ8fVpffUmdorglV4mW+TGRit/FD+/0176Qwy6yh55zJ/AEWGBMZ
U0ogbcqQhTzZf6//mCdNIHdAtX3FYl54hHPV2dXJYTDcvxsFVY2o2MsLzPj+P6QC
UMqXYZXfIJPoLHi7+bVmvHmhAypGLpgph8Lkl2vpe34uKO5+3L1NG9jKIoKk5BvC
4S3Wr/V8OZrkSlI22idNa3AEGEPn9ObDHw2qCYcq+OtTCIEjNbhq9RSRvy38FYXo
0WZVRi84aDczbqgKOZDkUZU1/QuURBXdAZf4LbGMh1ZQzf9xOCu/BJ0HV9bmY9Nl
aXxIFyafrMjBAtL4mzgE+QAZaF3gtuOVTShDG5J0mGSjg7tMywYZVM5HsyyTZbV6
C1oF/310DIDU65CfVPF71E7uoFHUTSgFap78aMrbUd5Vlw0uL3214agpKx4VlMzG
YQKfQXtpN9ljpHF0pFFiZEvEBfJZP3QeIgB0q0fb+FP4QIDf1iqKBXHnMUgR8KZ+
4OUcuXotHrGZ5B7dn77FtDpFXjDTB3Ltm4UN2FuPqrZEQFMsfWIdC3m8ToFhd0BY
Q0WKteRNfPMBZNqk27re8cyDuevnjS0IbCfoH/1Jn9MkMZsyFGNqSobynBAHIxlh
5oYgbkm0njMM/m43Rtd0etKOQRtXoFBE/1+NxFyfCQ7pcdu8DhYgWdnsu85Zqimv
SJV6Iob+nD6chPrBKd4d2C9HH3QCL5FxD+Syv9C/gpttvDMYKq+rs+dQ9cV58+kI
wPNzbxXe8HMGXmSZZZ+/PCZVMLxwnWMVFqg7lHsSRuKgPfFs3Gq/WA32UqLcJBP/
IQ5yii7knS9Uam+QvgwuJp+ahk2t53joslpGr6nK5plvfknqzf3QPfhJu8Mjplhb
zghVlSXPLNNzht8X0Gthcjr79o6Uylt18TEGV+EjaoEVBwevuXtyyRW5QotBnjvX
UkxVa5l7qbuZp16jIoOE7H8d6BDRneYYfc6sOsxV0WrHK3iBldaMj+rwtUHLvFXQ
RLHmPSVYZI+Ncd8tsy4bePut4CDQBDQU642+WtCHN5ve/Oz5vR48wbxJ+KOGsdfK
C46N3e7ZrojgtR7/VOQVkNwPtSSiJg6r2WQJxLtdgNlseE9NcTNL8w8fCIvtPzyg
x8ynscICEPQ1GDzWRIFbKnrzKBpNVfVADWXC3YhLbCORAxp/VJe6oai1MQaquc9F
WJ979t3Jcwu63kpIWBaa4bZ5l9XO2fvLmxpNOACV4VJGcP7ljiQJIyaAtQM6x0wQ
gXH5IUpO35g1/FTo4TR2hlcWrBN3RtcP/ZGQiF7crqEl3DE4UHUllNsGjnmQ7Y4g
OOtjnr1FFSa3iXHMcbIltJaC2fJYVTrYPSRTyjgDlbASR4/PtBJpTV1l2KN5RaoV
5w7RnIINVyotJmYbr6uL38SQuKOha3lhX/zTl2xu/yNTvaFlL1VyeZLoDT9PFyxP
FJR3KairHCLYsW0XBJYsTBp4D+a2xccGSc+JX+en49IRxOANdP8h53Xa5KZawsVj
0a2w2ZDgAefhMXOfZ8dxRONhue4N/X4BBV0LCGFGnewpQXqiLQymdJaEKsSU3bo2
xEkNdadNCnLNTN8ZnBJnYnllASrUMfGLLpx0kwoCkhMNmPyNf+QNVRTyCTs6XgjC
o0npZXQOSvEIprzWE7eCCdXu6TUeTeZmWWzKCUQch6+bO3G/GQx22g7T8hOn80L7
70n4U/xzFzMCTMSVxd/rIuhCaej7yjRi6lzuh59/EDQSsgQFBUWfZw4XM1jgAm2g
rL9b5Q4Vzkk02corFibaP5HBkRvwGYAsUMO0q/sROqzSZbU6wJqDzTjRq5vhTuLu
QFDo5j5zKH4mwBvcAYQGZtfXIG4/8Pe0FwWKrrTB9NeQe6kpxdkp4DbGZj+nIaU2
nR8iQxlxcIhFfc4MV+TU4LaeTJ0V9mZy3djtUcEplJebbhfhFC5GrULLvimA8TWl
zvbdqaW2Hl71OhPTyC0KR0RvM85Q8pxEmaUX9PWnw+lKhsLQSowvwGdfMl7/bcaa
FfTqKcIqN57JRoK2wC2SGI6PFIu4TA7GLndDIurIbTgN+wXS52C2dwAPNxibIsFa
sFQIuHc2cJMV4qYgsuInYMWimX6OYi12ttXasdEx2x1RMC5xCIj+Nm/NbyViGSaq
pnzgPEWWMyeoZ6NAbGacFGmlqSpVEaP0Y9bGKZj93nZAV88i2bF2mAKXgpiaFw+R
5Ye9g5yq6kVNJlNYWdpqM+65Bdh56JK/uCku6XSR5lrcHr/WzeXRnFnYxJSGNWfH
0xLlS4779++g28AzwgI/3ZHExIfEanbQrjQ0tHTuHh0IKQT7ZnvZ4e+VZxeJk6Pa
zaNf5dLmyGUtsRTCS6EMPZLQkKSSYawIUiw00ken3Jl5PbTiE+WzXP2cekM9Lt7H
XlspoO9GJoFfV+Z3g1z84eXJw0Z3LECkh8/D1gN2Fw8Ibyc/yWNBooufQgktef3W
C1raCZe6U0ZAjG+TJfLMOm2QBwuXhvsV1Kp4fXR260dGEi211MTMfsq/mM0bj0eX
xJP/bTTBIhQDQnGk0DdpAwF8GfAPtleOg4QgYz+UkcXhlKWmjmWDlGUm5tj9s/oB
cgxir4+fUubZxW8ZGOSZOvWnQcnb/tQBTGTNTTkFlICep5sBFqumODMNRugG5Lav
tBCHEYFJ/bKZ3hnPL9m6BiwgsfNAu1AhQyabY/dh4qQACE8apkNU2JMLLvngg6Zg
ZAtxQ1BjTucw5iS+97wDXzO4o28wiCqvUq4O3cXZxoqyKFeq4PoPPKA6D/GQRPsn
XhN9xG5Ni7dbEcE34XHoBs6SenIYlA+C+IhOfjemXIHrQyetvVYRY//NHJhMKdwQ
osI/tdWxiOsddzW5xhPFdDy6sngqpJZvVcElC10lSND+4w0Jx6RAFe356n3WggYV
IT+CRUHloYyuBV9hCJRzm34E3yfHRRyk6/Al7RzMTNoD+gJg3okKaK2/yv+w6QSW
Ak+pJGyJkKXo0YuaBeH3Ag84iI3zL8ct9nxYaRefsOKVUSDaEoMfOghWYzave6rq
6lWKJRoREp5ks5WcUgbBPXJn3Y7Ir24ZHz4wB35XH63jY1xYs+G5x6FKE0msuQ+U
uc2tjQ0s1v2vVt/YyND6hABs/BD2gejxE5UAIi7ZEteeFnzaVjwal8w1uoBaWxDv
RS0DYPdpYWBMlw6sMVp0PnEx2dnIT4IKZv9nsdOpa3AC9BwCDNMtjzVH2LJr1w2S
cw42caRuzjk5HGrQDQ5NTEkjfqifX8N4DW61wOjzJzifkpnopmWMFEZ1meIQQqyf
Tn3zvq/Qv+6weDtoaYTcCMJ8uDXna6vL9QCQAhOBMxxDAgUErrz4DH7RBVeMnCBk
vYDA2dRUL4n+OGvJdhTLgha1ShHK5g7seCgCD8DC6qRxXnDmyWV9mm2rpNJt/yFM
sbh0MSj3DWcF5TZzPaA5CXdRISmMu3Fw9kh7Ky2gvpPwIKUO7TFqu3NxeAuds8dm
IcNPrE+oyE0cskhK4w6uky9c43a4WIV2OamyqkGuDg0hysrGXVm+HbrMHD2pZrco
BhixeoL0p+keraF1KJ/lVERJrEzUiinByzEhSrFLhxBe8GcxB3RR6OF8MtuTn9aF
C2EU5cJuJalAoLPGSnFO7N3WdZQVFmE7/XN040+ZTzX2zrWP3YLL4XMW0yMrMAAp
qdUAh4skEx+HafqhMaEz/w7Lv2hqIIkSCzlamEJ4RL5uHLoILM8eJX4nRG6NpzrW
e9m23tcca7bBPu/oMcBLiWAVVhTwbKyQbRJQnVbacrt4925fu9/8RWbR/Z+/Atao
wgMEbkHr1VjXyUEuoldEGeKEGhDi2hccLHkWVE+2NtKLtGANHcNFsqyfuERTwLBh
rBJYKVjY4Dpo1Bx+8zTucybsXj0EcDJbvNT5R/9um7Q5rlu8nWcwEkaqLD2InqZv
A/8hc72staQjB2PObtxIfIP9tviLd9xAFYS+uXNyo3LAKnbbDgRleckQrfifxEk/
nSnV/9Mv0mLNfYopGE4SPcWyZptdG33Ozp5WLzFWzyto8jiHMWVoojVQPclo51Ee
VlBrj392P8uuWBV0NVIbbqdJkz0o4pTFhsPDs/SccY7ibb4gAQO97rOyEw6w+GxE
Wtju714ePa9SkQUrg8Nc3raqHUWT+rx/K77R/qkGGMQSdMylsTfAg2ILmDK8BK4b
qtA0lf54HAmSOUnvC3a+SPgKqeN8a8przCuKf8wW2XxgbCIuaWVKI9C9YT8JcaJd
9aKieXo+9O+7mRMt7Gdp91RQz3oS7ywHnTdpFcBoaJtKBOQAs/CuAQarK4WD2fLg
ZINy3eAnRHXZAmkT16hc+/L6pZ8gXsCPVANmjaN7XeuzmRr6G7e0aPBSOTsndF/3
i06V2MBY0j+MQX5EgubNsVi7zyt+f7FWuMucmFFZBt/HOOm14lH0ZdPZoWwRJRZB
HoQ7/jQC2uocDn3H5f6oWd0ubwhlNowyucAv+3jSXYA/AV83DWiE09NENZwE3hc9
V9oOrOPbif7pmIR7QOP/wp60lg8JuxpiffCzrC6c/ETc4SCBpOgtPNRsBW0Ocm6H
HZEbvcxARzDmJbBL2xBTVzE9zrWLSX8fFREN6rMIF89+WepwVHpNo8msvRcKEz62
uAhjPdfnzlMhB3gB2oHEHhBsE/vmE2dESqDuD7xqy2/YHUggV7Jvn9C+ydadb746
LEAVhxWy6B5SgiYml9ZFVAh/eAGN0xIy5nclzj+vKvUcQeaHvwLyNohtMzuzvBVh
KR0pt5IBsSL3xaW1ilkBJ9y2bw/skdkPQLbCLQrWD6mJhqXI4jDkN2zEw1bz1nBj
RTlvc9Itv9RO/i2gEXcuMWsXN3J2QABwZPehKFBnovouyVT5HaTa4Q5EI9Lg2yG2
m9IbJd46Gruv+At8gb4PdoFUxpTJFa7BXb7u46aZ8eSclzojFeRoKwL4BSiHSUaa
S9NDgrFVTwrT9fZDMRZOmtfN8ZKC0M7GzoT/JWcvTss8dQxLzoiiyjqi1+9IgMC5
4lhgJKv0XIaSB7ZC6F2bJxsS/NAm1REi1ECDFZSuwmOcQNQzTgTfonjaY+wBuxcz
N6tYPP/SObtJhMeCwLsaz1IVvlcxoMUXTYovDEuKv/XTtpQmR1z5CasvZGehhnpV
VQhcjniodT8uRNsnKezFqm506N/PuTvNno6zisFldzsnSSJQ38Sx11vic/Pk7HJ+
NjPnNEII0wsO1KpfleHa1CUrxHTfNnDM0VaF1PLQeWD0zYslbByGstFnu8CBIj7h
pcUkjMXV1wiehaEWXIMJQp7x+SYVz3NEvFh+av2xKFI2kHN0AuQCzdvnGWekRcTk
fDlFkQRzrvVLNKdLYs1S5R79JRcxUW1pxHct+aFA7/ok+MmpitFegHi97Kj8C0+h
JbarhHrhmhXQ7azSYMIRT8kGLDzBeGK+1F9jhAy3+7C6BnWH5vW0+x2Jn6Hpewgv
xOk+kZGsgf77QnOOvvfPAV1ihrDfyDIzpICrbZ1nlbPn38TWkjl6u2RJO+iZqNg8
4ctvjr+2+bQcnNBiqbi66g8Bh2QTiW9NuFQ9AvPxl3nerlnHZjeTzHijfuZ74WQS
pRLXKtZp4CfkgghdCkJCk+H1oq1kG4QkheJt68SAenQaHQNdEZq7f2Pfn1n1mapY
zEx7GZU2H3vLBKdju6v5HWCUh/7vDnEtKAibZ8DH89P0jajDSTHmbDwHaRlTYXuz
U3HPItaSIxcNWQzdFkWhhhIqcUBubmONDXteGnSlxiXsgI35aea938wRNBGdtXzj
zqBqQ9AdkXxY37KiltrYqhJ3Ay1lKiA84q1+lk8vLPKjC1P2s3TxOL8xzbZJ+nJ9
jyO8GqsJF1l1rldvUiPrmJ98nEoH098Vj6PRBaRKz1n07VKWnlMTWKDhvtc8tDkI
ZsI8LHmzRa+pHWNtmH55O+g8CsPKPDfR1CjnY59dx25q3hZPSZpbXoToasXiWMlu
qBoyFIZOuA/ZaOm/K/zhRVDXgVZE8cCfUBjb/qmSTLwvjNm5ejY52hFEERLuErp+
OQwqoiwCUeImFFy7KJm9O7wyLi/knXUTHD4Yr5SYZbL/x3f2g8nNgrkHQaHsiPmg
wYm9zcI7LKlAJ3okpp/z31dJb3TMUYivVrC3nu1lYYq+Iqz0NYjkQluYqIHejlFh
rJLnXC3ZislhI6pEhfkeMMvR83kFy38vDVhKhUfPzXf9zu7h+Wj7VcbNmBfnBFA1
205TrMCbKjUnTMww1EvRzCPHk9mSKP0ohsci1s6dDB3vETlOzXX5XRY5SkstQ3iV
3KSZq5cp8PFJNvjzu9I846R6xX5p1NJsQ2703uuuXVx5Xz6/hbZ05KyWLJWoh19a
4tqplOEEJ0dq8eHCnmISbCGT1LzeK6kVuVR5GA88+E3L9l1/ZOtWI/9FBSdhRiyx
efH/6kkZC2QeeqHH3/e1zYSJhn2D7fXb3YeBGxK59ZcZv3eY7YCQyrTSDiDEstri
CEE9NTcbfYMN+mmQxPybf93CK61Ql9NCYrtj3n8VfH13fB5p45+dVrOh998z0cA6
f3at5wXeJKdaORN5ix+U+VUkV93D2xSEOxQQiPNxOOJENOYZHM9OI1cDMEmnPb3Z
1LEXabRiPzFRy6MNX2FfUfiZbkPm+sVjdQ4D/b9Uua6Oq/v10oUxxYU/0YkenH52
Ib7xyiSynTMvAa/05/WF2+KJRXARtKp+e9XEYHwcBqIM53mpeOW4ErJwoulL1Ms+
0KEo2HtZvi3JfboZB/fyseXZLsjcFvUPGPhxWPbV7L00qpLXRgjfXBSZQOdf91vi
JhrBRbgWZ2e5juwwLVVLcWwsVHlN/Ts7MSMfvDhOhjHCiPBtUdkBSs/WD8uKy66e
UrMqWw7cDJfZ+fpmSe04+eqd3cFdrN0/ZGUWXywExIixv4uM+ZrDJbYMPB+yAqWS
6rfKrWJgnwhx/KQI4jp4qSqHAwMJ1xqnFSYwWmPs3LUFk+rFcQX42QaqjbQN8CXx
br910Ots6087gZJTugW+qrexSF93thD0QiqTxeWJ68O6n0hw/YTqVY63LS/Y2Bjf
CqpZrA2r3Y4E00SdRXxg3GPfS+HHfERKqbXXdFs1PJehx+kpvM4lRWyRoUeJZrj2
i51yktBf5fbHYLm7PLWgK6oyK2Gg4alsNPss4mfSqC4iAc5Wuy7b+/XZOuq+OFkf
ZNhPrtpuVt2rqUAmkyxAwp9Ky04ll5Rn/+6DtZNLL7A/tQKXvK2bV9dLhDJGpKqU
7afxIaqS2OJWI1IAfcv0RIyNZLIDGXPTnFgqwkI89OCgWGJdrFa83oKwOAi4dPEr
hN1TDhfMMDNziZoh8xV2HQBsX71uiPhVxjlqScpBiaQv/RawLAu6E2Erss7kstOY
nvnpWjirDnjElGIquSxbbhF6S03Pt3oRfiOqAkfhuCaLOO5ODVHjAlcYGlLXtZEq
KyDzaCShUHmV+nPnIrIWM3uYL928WASccIWJNbq3aOIHVHBYQUIwU6xDa4ukpjGN
4W5jZT/Ar2wsYvlcNyKENwqHdRk8wrrEXmalFo4ryNGYn+ep7LnJ+wAR28U1dZD6
NMT9ANQqRM0CplDMegh6LliYqxBONwFzjVZYssaMA57rzghiMgpvRtcu5SjZt663
RuVhe3dXGVbr9yB/E/2QWZ7Xo7a9326VOuXqqcLtSc5QHWpJJYVx3UHESxXK5ihB
eIOkEj1EwLCzsllsFPBZBtZcJT+nVVkuMR0f/7BN8ZKWLJwrU770aGZFMmCQtx+1
M4xTDMqMZ1p7BYk4phi6pOVbjRLI4LvWJKrJ+JzOs7I5rCUkjSrw2b0FKwBXKcK+
pbn6ubRR0IWhA/VKVLUW0/O8J/4AEiaEqQMqA55kv+IyZF5LsLeA5P9bnzAqohj+
djKxzkP+pp8N9+sP0/UyBlQwqEDM2uu8ndO2J0u9+qAFVIL/EmIfR0LdeLhK1rjg
XBEKI3cV+tY993MOHN8pdWhpqgy/j/i3jGpSv7vt43eg3P0vBzscHjJky8SmDd1t
R95XzsnTA+0l2f6wN/bOgsSg2Lhuwp/O9ex9dMaymTld+2IQvPsbzPcoH2vXyS22
RGiTFkgzSMNU47MaCylKKYJu/JrKVakCxOv4l6IjWaUFyibmtNy68/r8uFd8W0jk
ARdD+yP/0QpoOmi5Y4KajmrwQAoi+iHGNCdpwIAbm8PpVaR3JrFAalZa8Zibgvue
zYskyt0/0sOOFvP2u1R0rdN5oxVifRfk39e6t1h+L4QeYUD5Io94MCdTJP+RtUqo
WJFn1UPMU+wQSjS+nlQb1+nQpsajWdOXeseQEqkOlCMFcEwiNCdTPkCKJmWvyxIV
oE/R1WHR8+GdKLAOWpYhKE3xLqIQVrAEwerVi7fVxD6PcXrg7zV5RU8BLGevLfS6
ZwVDA/2SQ1U3vZFYnsFDcit/efl4XaY2BLr90ANzAhGg2Q1xufyBjocBkXIR4guI
7I6IZC0DF65Y5Wihdv20PepMs8o46aIkXPiE+jxJ35gyoHJhv1vTfIBxVKMR5MbK
4I8rFdMDaTDjxKU8Xa5VS1pn6nK3rg7t95oTTLmsia3JyEcvRsV1qXCwWzDQkEVq
HOOnpvbvuwDIBhjqvjqWnSa/UK3cqXu6JcXWnLXVpfARcv/iLpSuUv/sh0fa7g1K
r1OdI4MJ+P6TFRQZpe1ytW8jeZ0co1GeBlWTxvdF6JqoOm0ViJp7E3f2KLQIJ7c6
/JYpMnjwQLj1QLQiY7BxiCnt59UMdh4UBU7e+W9TPdNy38x/LiCROxZnlfJttWUt
ko22VPrKoWhTrT+geF8rTu+blR9GXU19bA4I3RYaG3J806UMdN1DM8diYrkfi+iz
boAEnMPWVcWSCMROs2P1EP0925dZUJO9mH14EMZp+yWKi83GCCyZHTdMga8ieI1j
+k782y6hqO2FjAkQmz6zTc72U6Kzb5nG7RxL/wiye/gIatZJzBtXTJ/PKDXuq0HS
lID9SkXiEjU5C/VLzlVk4JLrb1mItFinWkpVq4Vi+jtkNsuEYTHioJ0/qOd/PkyM
rYygy3THjrLEGWzYdHUYBw767GFU7spHY08X1O8d34XCvXVpXvD22Ksp8j12/SqP
Bn76N3PJGR2WQOBcibeJ+bWGzI5EQadZiHWiHvAk7mNwP9ZLZE4tQsx9fPD35aBm
7U9Z8c/OedddrEU/zxLhIUdSAR0RXn41mWw5VLGQHRGf0awZHSPRhNBijM1q+CHu
m+7fK0I4JFFCSiHi9LhokzusWLpOC+zfl74g0Dfm/BUcd2Uo161hbmzpnYQoEuPq
WmGiRRNgQOC9GT33ufEoHH0IeU/EZ5WF5CphNS/cDFh06aKwtNAvwlMsN9Xt+xDy
gK8aE9qc9aQguIf8xMQN+jU+EMmPBpUYcKoTs46ef4lpm1LTR0yep6Qe8/0XBc9t
udWCPUxEPdKaVa/YV2yA3zUde5yz8V4g0CQACAFAxfL3FHqQvhEnWmR7kbAQ8Ovz
cwayq6s+q27JZvnnyaPgnQ+IsjxZi8T+Zw6LHBeChCrSnwhAVcZ1FS9tsPgz21aO
rKu+/+sXS78u/7B5CNjKHrsyhRMoiqvrJKJ8KomQRTInd6EBVLs3iFUBKPY4jVUo
/qfHtlboRtyFQq21zMSrPEeeBbRH/6UClCZbWAlCsNwEgk4D7Pob2T4ZFOso5Enj
9v8l6zOxD7ekikOeJaDYLt7jZrVsD5AQdUCBk5Zk/pxdZ9LnidrOStuZiy6onF3C
hAxhPXqP4IYNsIlG2jGr75GeDhOJc96yko6XslxfTftwDc1ZHozZ1QWQ9oxNtZWF
4BZvF72wY9pA2D2RbjPcjw2cwKUYE+11reo68mRn5+vn2akwRCNzYoaU3X8WOoio
r2pJIwWGxfI0GdalD8teIUMGgG22whTJ7l9wow1J6XD7SfzK9IlWh/ZXaEVZ6Gro
P1ZsHIolySHx9OjSsyo0LW02HzjQXtVxFpNnypNLcUMx+UMoRDhGmmRFtC9m3OR0
Y+Q82IcGd1CfPBPhraXaiqrHyKANtvMffYt+3Jud9uVsvyreOOykzjCszNn4gbby
LfJwAeFemTzyIZ2IoaL+hzaG9oRUpSlCyyufevUJpoGxNe+5Mzbh9TPVlSfnJ/Cn
+FSd8SebnKK1fpMI0c8iOS8Pw9Mf+GGc/UFzkDs7xOyPb04ErG6tjtUFVepywyYY
Hp/ZWNhC1zdqPStXIGe1tSH1pxzt3iHVDzmDKo76JFqeYTX/ub9VKw7nJDcNAUU6
ZBIxbWV/FsDVbQPlFwDaIy/NVDiCK76guSPoGdWKgnalHrRazukSDyEKMaXBxQ3y
iCN7AaF7Z4SA3qFJ784Ud9ILDc0uniKivd490qdAJgRxqdbcUmuPbba/yX/5gv+d
KnR7cWm1OPIXLoFvxFQoffCthJSYhcAQt057vOSHOnme2o9bC3VBKbLkvvyMrVlH
uhHEyEnnIhavZXSUbatoTJQGameTomZBfHUXWSC1DQ5rMQceNIsP59gZxl5Rcm6c
xM2QTckbairFQr/SgSRQiOpDnKdAadapZjnKmh2CBuVtxsR6FSWnqoytomIku1M1
YNVtowckIkRO/0rcsTKQITbEfPgQTtwLix7w2lAu330ee8xxooac0ZmbO5RF8N0k
Dj+l447Kb9rmao6YhRf3vJHVy7w7DiVBFiyIHYSaUus/OPjYv5ek3/l6knezmatQ
rgRVE0EIR8z2rmLNju9GlnhU0IRZUR1+GS5dRrOgHMvT9WduIpk1eb2l0R1abiWe
mR5mOZfYnjx8JVklJ7GtDr6DwVOmbYXZHX4nqpVMBQBuhD2UcGg3S1tSp/Fv842X
mZiSIqeSoRCQ03x1WY6tEzWBgJUj0/TEtcbeT2VEDamr2+4qD9pGhv/WEL/SGLdE
JQ9kZDxietQOYep7NFXRPK8iU7HCnB1R/E/11AaV3u8kWF6VLPwZz98WMGGquvpa
MrqHZQGxxvOUUV9wptxpCsFM6pM7PMeVqfb60BJ3BwMONNx4rerfJLJieI3R4mM1
nAjp/R5+d6PMdIXm+Hb2/sILxm7EyjMBJPsDba+uxRUyBJrcDfEGoQ2GI7eydt7S
d1Gi3/HSjqNznHrUHRGDak8FXHLdGDE4XnlHJepVTZKCQczIomrNF04dWEo5dz38
d7aWkyJb0Kpr/xZa31KnRMkNEfXZMsJpv/a71829TxWL/ax8IplAU4kklHRqk3CE
CKqqiEdxqm3l4IC0z/Uzinq/KFsEUqPRPhWsI95pBfymCS9v6u385zf7ku/0CTyq
AFeUyvrsR8qyoktUyuW6UXF6xegyyTiY8NtyyRVRdzFsTISXNq7os3crt2/0yejB
ZWeB0Z2cH9zbiNSuOqg/7pCk4088ommvm/tEAqUqQswGtgpjzFeEQk1qXb9ZvrTc
g8s0imb4tUUhvafsPzAirZ+/tpMJZzztaYV2BZT+JXfkmKq+NDjcKYMiU+UfU47q
UedEym9BgosJwNkrwh9c4I761eiSjcpjiTLqkE0W0cWJll5qnJ1kG1qlWcTs3llL
kAEUzqpo6SJOxfqKLhnNuTh9UGKxxbHa9kYHwORgz+5Y7ZUMbdr+IUBWuE5edndZ
RhVRp0XD5SuyMewPjBF6kIKQuT8U/sg+EECYPH0WvgLe3sSTZo6vtNaW5XnPMLsG
GYfFwC+9IsrIOatrUuStosmCdUCLOucXwZEdzbiXqAnYQs1u0okiqOjTYz3ERLIS
EsROaa15yioEje5QYpYwtvwiq2/k3Csjzcqo9Y2iLIOw+KWIshRWsh2Cy3sQ8fXN
NFQ0GJcVNVaT3ygmTp27NZIB2psspuUTsUQ1E4CQjazmBuAvta+Pbc0FQ2YwVy6t
iVE0ya7EHX6/Fj3QJHHB8PhAi2/8Acf4svCiZHpxOWJne6IjVEdYYeQQ4SNcZsrG
L+eZ61v9nkgmzD9kOTkhwISz7iFniDV6uhIiKoRXrpbQLfBFvOxg/RcAEPGPQwa+
twL3Wnq4Oz7snG7O1iWVOyGMYh9W3W6KBAHCoG/in6hKg5dJvX1PnPF6+3DN2Fpq
Y9zhP5zdL3yjphDuZHXx+IdYId8PqgJVj/aMwexNvsQw/ywb9bhwo4RIJhXn2kc4
P4sPYwjnsQTH/j8opAekMM4cAuWWhyz8Zjo2mAA1ndh2wcnW+pQeCeNftEPmi3Ha
vgRAAeoaw7b8xSnNvyivrnjrgPD0FlSf98byLc98HddIi//cIJjB8ju72t6oZXv7
EnafT+K75HzQMSB8es47oF8v10/gB4AQvRna6sxHdd/q4VzrY7c+JlyFviKxKWhq
+Cn5a7B6oznsz15AlF7e53Qj691rQPTHBe5mEt34XUp2SVDYN8d3YVFEfdgyJWXi
DInlV4Nvx2prb1d5dzQrf2sAMwP9sgoVm8RqaPYY35AFV4W3x9p7/6JqrIxpioEQ
sPPJA9MOdm92Bh+PJlaW58uPDystZneY8WoU00HegeRIRCnK2eSXQLXhqOtM/my/
qUKJHAXnY2P3SwgjyCFdBKQYVlRhqELUdMcRDUDwEE2r6/kUkk39VxQ2CjLxVi/0
U6DkB640xs0bwWHDUm9zYyc13wEkLXG0/zKdYkyEcR1usVXpeUPrWK9jgSNK+9L/
WaRslghBK4/F6QnKa2RYyY5RvxejHkldR8gbg3Ttdsxm0yP3Iz6y6jyUQTRgpBbI
t4VOAem3mA55mZ8+gfFZLiAfq/e/F4yLOXkqITqt/SwhuwztB39EsiyyC+DiGL93
70VyEqBnRxIqvAZewjwZHRPSnhAyY9xbHAzJi983yx5g+SerzYXmhOXO4JB3MlDG
+3YDWFHqIIIEDEDLA1g95cH556CKecasivj3M6jGfILxnU9tBjAzeL3xypdrGk66
HN0M/rg7nTxx7AQTLMs1ZbZ01YaKFa8E2Sp10PxoYWy9oumsLzgonIcoWHMrWyVp
JEKq0UwjXHWJX7WMwhwY+WsEkilgShUZHqfs3Gwu4TTD0XBoGvkKaHzIzHEg4gic
+qs/lCOOSRkmjfB167GGDouWmgXuD8VLRzDlFnrO8HGqCDJ3im5vUUKUg2u3WJb3
opCVZXRl3/xT5oFq1Bszs3jYRpN2AsOPaMCBL7ekQz4GlI6wm9LljFisbW5pjONv
NCUfHLIS+HA6XoS+ZNmnIu+UgPxTwi9hD9YAxbQqoPT2YrNiZue/HByzsOa2coYP
J2IE14bwLD1K5JYJMD1JwIsk77JJKq3z0kCTKOaRi+DI6Jw2RdP7wZceETWsvyse
kTxXc1YkNouo+82PDCuc9ty4xd+pL/VT5AVgFi2fqloXi+kwip7yqBXnIGbzfZ95
zlBWaFFE5JY+FsrKVgv1UHZiNWS2z0ACYGz10rWvEuN+tpJWyHQ/CqhOWl6LOnog
Tv4jyKIybJnzMysdfzTJp/s0z3xqyoDdfoJwCrpIlBDs+zA1lEYYTBoaAullIKeP
gliKRDgseuA1N2/7fJxkCQ+/NyJ3woby41td8/49c2EEWqANRgDHXW4l2w/SXu2F
jU1zieshCGqnnlFOkveEfx6vHJu74E3Q7Fcd/hLLr2qdinsW46d22jew7JwnL3K5
7c1+s+QpbzE7khL1S8EQVKNA484lO8XmHMcLDs8eXC50mEfc5lVWXnCV97yocFUI
wylXYPWZMzFJ+ttKFR5bhwuxCT+mwK/AdHX1GhdURLfu2yQorBco/FsSeLPzHyg5
C2qvYpmsUW3IDNMThpk1SUahkvlxaFC14kmrftfWdv0SFhq/49xu8BNy913LwzkN
uwzZWdbuzqUQxkZ6sKrlFhmC1ojXgZC2RjzBA576WOYwUrdBjac+2+iaWV4dKnrF
8eh5bI7NGh8Iz2Lmy+p3G65VTuct6LE2bSjN1C0ml8LHr8VbZWjSR6FurPhNpld+
PIJ+RhlmJkgdTvmXPSy5GO6jclpcvkGGNL22N6Q81m0/Lhs24Ym398/Of92odFkD
j7U/+I4A4sKfsbdxrJlKVlZZd7YiN8Aud5SYjNmL/iMQbOABorOMT2/AYV+ehZLY
dHiDfzwo6yVXTvm1hNgj8eXMdPAvaUcDVQaOGOGr1aTZev08OKP5vCg6AvjlJgYm
w+g8ZRzFI36xmD3yWKX1rkDLsXG7eh+SlHgkjvKLIL2SoHJixsDAYDiUMg0/y3l+
F1XphUISP+JLpUkhpvOxDOhYdrQKUg6S4IVabAat9ZLvKa5Xu710YM2Kzv7aju1k
8y/SopnGgrv68BKJnuNYghVp8+YUF8qeYnvISyM0esvBdNHkVsVTk4YrWwEzsO8B
2T2MsDoM0y/VyN5v6Y5XjDOANbSYYiJmmudRyql/BQ4ZdodT0D/guBeYcC6wOBm9
Trwsh54oQazHZzGVNKoqA+9HDXoFqLQiDbH/Cke2ZeWX2X5mUcHPX1tYPc0WXsxR
f2vMfLhDGxPDDG5Q0WSeZmuukayGt+dWZKlMkY47ZUfPwzdI66DOsB6xIPwk0qQR
aLDgCa8ELQu/7HqnYvYj/X8vV18t31+dyq4fScPJJZXDjcCy0NV0UiwkMSq5Npyg
5B3yZSkNESjV6VTDXyK/VGNLP6dmXKYh8x5U5PaPxJtkZFHgR/8ofRKSDiUwHjjy
bffZOnhzJfnTljwTHsNUhNfUdEDQUr2v165FuNRzH8vJw6+lqIviPftEBh6XqNhp
6zJZuxK08ijpJlO5T8Rz0q5Qui8pjd/Qx06HiNRF3vHWZKCjKHggd4eBUbqN8szv
xoM+Way5MLBdmnl9Mjo+PHUoRUERE5blPRiZQtKnKkFgq7QOF49krQY7I9BpfMSr
5R/UOIU1SDMz2G4FC2Vq9C5VR+MZut8a9CjMXaKHqDBqzeIAXdeszB3rXhx/7A5/
j+H5Nwo9KmS5NWyuRyfPe1K//0W71mbuMZtJFYfBg+9mHajxJfnr7HzZ+3hYOk4+
6szOBjOYnK8wtq+agZyGhYNsY6mGpNNCpkpUke01sG5kp0Xd0APbQxVkgtaAiHWG
NR7oBadot0+5VBMoe2jZ1Dglja7/Ss9zhR7B3O/mdBUxyA+W2XQiw8Uy/H1T7E7u
iVTWNqZcwnKCsfS1atdgneicBhevptnECwsYh0f3op97/H5DrsjDFj7PFMo03BTo
1EDP49Nh8RXK1uXCbJ9debOBhT7HLSS3RQsMRYCGEbvz0i8HaBHzl16IxQrmxbDG
hqYFw9D72Y5m5OZixPS1fYpItAcCf6izYv9zv26S4zZ1fqbByIxHmkQ6lE9CUvbn
P8Rq2/mofNJs1pbskBRZKasi7P5A5kC8VcknzCWhG8OHdIWp8BpYRfOHnXyMlL+T
llt8MH/SXhzQbp4Qqn+JYoQvkuYY8ODcizwud2fZfPfU58gQ7lARYG8Fppli7WIY
GKDr4H4xFf8/6Pr5gLCDO7ntVvk1Q6b2Y664OXNNd3Rv80gvsj7zSknqH0zglP2P
FLJWUaDTsqYDv09ncpk3jyvtbrnUVHpnX6v0PgeES1rs8E/aY+dOeWC4TcIfwA9t
fEyYYeQPf1q2yViU3adkcjNHCjKkVVjrIBudFBZwa3iIWVgRXPRQlqn4FE9i5Iy+
gDX0WrfvDtMSxDSNl0MLekAsEdmoFmsdECtu4G3COESFmEUKEtyMFnCUYOYSG72y
gPbEh6H0KFaT1+WxF8VmHZl0VdOklPoHxumbGswXK7KlEkDN7UqXjBp2+veU+UIi
9+720Td/JCDqIJKMJAEzHNrDeIxc+q4GdGi9JtWzoCHCpPJn2yBPKjf26PyLeWAD
0tahgqgT4c8+HcqwJbZ1OvnGUZPESBnf2M5WF6DgmjAlvU9TMhcSPaFihsVi6WwY
9x0Cbzw/KbAhcjoxPj4bwz5KU/MAyz3Ghap429KHwnrXspPcTP41mCUUaRZFil/H
KJhCx5BD7AnPZyb3ZEMnpo/HZdMbYWuUshcRPJ7tvDYRcbu20lb1ZnLNwhDFkZPC
bfPd3ENNnctpxZxpuhmOSDOrNkBFqfZbI2Nk3XITKTcg6oGbwPqyDerT127u7Fgf
7ateZa9JGMHOIRstqxi2Rk7Y8rbSs+83VzUWPRepzSoHsO3kYRj9LeIumvJNU6bj
T2P1Kx2mhzEQIxYVDzJacZAIYYHHcGX6PBh7sOOrxoTqCEkT0E3kt1jtGEAzJC8n
rhp4qFyiNK6ivQbf9b0/44DP7O05xM+rJ4lP23Ukq9bWmwkvMDXOqGNRo4VY/f2H
jgH52yXrd7FcZaaswiFlSLnKMzbdqMUqJTAPDt/rgq+ClLM12xqcJb4zqFApYbOX
WOGKK/xRbYZlIqLcaafOMrrCe8eGmNkb6LP1VvF4gaFK4IFGWhXKkDqbPTEu19oL
vmm83HhhLyafiWnqZ0z6UsJFQRqfMAsGu/AUOtS4ChkRT1omwU/afrhqgfUbGxD4
WJOTq9Y+da+QRIeR31KpwYREBFJw94qxWDrP0kM4nrK+ncDQMKQ33iQ1ldiFtfl4
nj5mQLANELt6yTMqnyVDOBcQx1ItgdtEEU7OqpRZq3T/Ha7l9JllgaoP+SUb2hi0
J7aEF9O6lLicvgkVv7kTgofLMMVu7d/HlXcLiieqDheN3BTFJ3juwAqspPofrpcG
c0BavgaAkk+xz5p/UIxi/MKlyJMOXtOIjz+YQBA1rclTCgoCKlsMELzfbgaxFs6f
/ZldZ8Q8KNIMalwNzgnZUOeY2hE9e16iZVv0YeU1vi9z1N0HxX4dCqpreDkT1b7Q
a5XqVYlHk8CKOI9pj8owGd2EgjNgvIo4GsKnHt239S/URu0Ju9vT81v+SAVNyHHY
iUvo+9CGYQlX1jGZ8YFO/3ukuuhq/o67Va26aAMdEQHjnZ62rtYpwXUJmzLIA3sq
CGt/DjpJlS/plZRi2/wp8k0XUZqg7WSH9HYyKY0/5bRtn7t25D/acRNgS5qwh8HQ
N9MBuR1eLfOfIXD6Es+AFaaBtW6y6s5BuOUw1F3EyEk4de8wDznXWoLMwpK77ZE9
ZK/W7b/iojFNOerbKwkmL2/c5JiSVG6G6ji9U9ECnQc/SEBqbG9RLcMlBPwSKrB8
r/Hny7ApniIah97bX2DZI1QqvOjJ+UxjnwqV3PRw2jN+ygk1Mix1wa9q/sHO0h6Y
dM71dxwKtJVctsuUQS/rKUWos0IxsH9lkBeGjTnVT46skmq0wFsP+/xFfhRfsMZn
Hk78zSH9L9CALjvoe1y/EsYshCznb5h3J+J4rIcS5pS4h4/ErHTB6mcUebCRet95
J4EDOD+d36ucNFWgkLcVG89QvSONKfj74hMXAU/syfjhtiZA554p5JHkW+woI2Hi
wpxUqVHm/owl39DXsYX7OiWCIQUsk+fv+4ZNUPPEdqHDeFzAFouZ96ozAO8WQ61b
nMg+HM5YTR8t0fW11WxZSxNui53A+wZGWOFvMGQBN25aGFkjNqAc3b1kb8Iz/q1D
Dg7driPw/ds4+F3fLVOsbRSJ2o7/VK8V10YDSPMm/j2Glbl45w+am5um08blJCR7
jjiq41bGzT+NoEpTJOJrpuWTUBd//eudAJdhe1AAvt3YrROqxoYVzdap2cdkxoSY
I51wit4PJelXou3WCHl/N+s4U9ce9yZQJ5X+qwvyDXhmcEXym5o9FDi3kckkbYwL
P2aCW0L4PfRjblk+Rau9Jb7UR7dtScCZqWWtZ3xFBSM6MrrKwu+pCTcxGf1QDmEv
xqcUesc6X9LcvP1WS8kv+/nljFTCILYqumEuAilpKrEfqpLPEUhMNhekewQ+jNkc
j0mVBCsJX2jmly6ruADbynSyaXcFunBN0EKbYgl1wQ47GaIDokHjeRTw4tn41jsP
/zVknUw8SHvdyLqfmMXEbBTWD8LcEQD2+hLy97B5RIDQs2Ioapq6rcQOwMdoVJ0W
5/gmb/BgxUQ8a0ITah+ovsCgGzYu3fMMSN2h0UlSeVjLNiuts58mWsdC5QIitQyP
gASueAQJtS8Xi0SOVwbKPlwJXok4n4Gq6oFxYKJH//pjUmlOYFOioGXNYpqYKsjB
R+kCPdurilRY2T0s4xS2toU4Zvq+dam6VJorlqs5PQcwFTlm7c5oPV+K7LorSyLp
Z4i5lo7b1gZlo0hImcEHonkiXqrNm7Evc+UA+JO+aubeGT5pq7vm+k/92+uYzd8O
eZqj/L99kiUXCFkDUnwIPZco0I7yvJAskqZthp7vWEwe5PQpWhukhlf0+N7pa4Ml
kTNPsDmSxpQo2sHC3h9SIL2utjGOykqS97bXBnQo4EUJBr/pBwyGMeN50Zfr9RvG
wCoDXxLeTI/5IHgFmrnXollprdqDoGS73wwzJCIuEtZIP1RwfrOQmBdjJ89RZDs4
tvFs6gtfEtwZMdoFjrTcPGm/aBBa+tbIu3Ur0odnx5pTmoZ5RLvrzF5QvoqW82G3
OvuE44C+iyCWBShMUqR70bGdDBHv/XZiN1KFr0lT9HNiEjh22WY/rS2ol9bntsd7
aJfOLFplZRZ+iR/NLzXqBPfdg3uZ7+7eQ7a+fqr87JhmCujOrQY7oZdKinQj/dKk
yUO6gTxoO5PU4N/v05Z8O2gaG6b3IdzIDWumJWNFjEceUtRsToTm/ocwJJx6UGeG
RmifXun1+pF6nyRJY8pj32uyNTovEphNzjcSozFHTWhy7pgt0Odt9+zneUjKDY/F
nCXrKas0r5flYzqhlR6G0M8T7UAHJsfq9gdx8asrvil+QLqVQ/ogE/5aYkpCxiMk
Z9POLXN3pik7JbQr3b7oRT1JsDHgd9D1xXSJjNxB55X3zf+PNX80tM3gr1ZTRu8k
3yH9YCKHtlM1VzutiMPflG2rxOZUQTLnCZWr5qr+NfEqS4lRIostalC6VBC0iDWj
QwemJ6XExiztHX/4GHdbo0Snybzaz+zGwJxQoeXH51mn3UpgRjRicn4BeF4c4fUr
/Tb+4KJQ2Hb8Ljd09M02oCCeSbWWeyeZNck2Hu38OHVk89bl8+IyLsUwS/Hhn01+
vFnP3xLJnwmERXEu21tHJ+fxva0wqY0FZDz9aoHrrQniu6m7yNftOqs9tg4Ei3+Y
EdaVLjphwTyJ/stTbK9AR2yLAD9i9yYcZDxTUs8DUv4/v02Xtz9tzKNPVMnWCfx5
gmp752LjHo2Y3i7X0COBOWlQpHe1wIwdH6ZFzmNR0+jY1OqMmftE66/GaYiJG9bl
CJzbJ95sC1ubWEQFz42k54R6OGwvzAuzA7dYgbAikxjUdGcaegwSWUkYK16WTt0f
KfsB8p+pAgAicUnWaRJscvxUkBKCk4YiTytKVSH9K08dMhZsgmOuCVB5etY1byiW
yTeat2kjYgkM++qWiGKhfQj82m4M0Vx0Ml+82Q1wKKeZkoZCIW0QTe70BbwBsQuu
dEA/Fk4+JMxMY12EidTdtTURcmK0ewTGT0UAwjSG+zOaLxevQjnIfnqaY3QZ/5HS
JMzQs26P5JCIhdj+AZvCD4oLY5XGwZLwJv4mWRDskBlXZsz8wfkiJSU8mTOvyzcr
nflGCu+njowJi/QUE6wI7/1Er7Fr7ODMQ9cPs1Yn80nf34SB8HKtNo1coG4nHGsG
l+QDiTn8W88OrJP87yTVIpA6oNio/2rIwmLTZHo2OE3CxQPwKYB4AomRO2Qv0/cT
2Rs0jnugvwQl7zoFMjwXxTdKGMJJILB21TYBN01nTirrwsIw+ZdoPPXBtbsW1TgC
ZjXMKhes/wvBU629EOMs7PQo3AG+G+dL7aKxdcfdY3xZ8fqVlStVuwYH0LKLoHoG
VcwfJggX3dJWw6vNmx3c8IbHVyvORXaNCgYtazNXAwnOv3pgpN2j0ET4ORsoTMM2
3ErhINztZ6MV4730d16PnokQrJ7+u0KhOQG/FrGMdVDMYb73znael1niMWa1CBZe
C50E4W+nlAMk0PFcJYdKVoYlRIpf7rpRrKBJcU0BhRtOCHGkMwvkS2iLl6Kyyr9Q
i+BYT4gfbIfwcU+IuwZDXHf93idkJe3yjsWnz4rnixWjX9k/IPzx9h2+RIsqPhDm
+pUAQARNoebuPr0i/ege/rTPEMM3+asY/4AhO0rVEYTvQTEh8jM5j0FiGPOAXdk4
Z2aHSY+FrZNcrX4pJNTmEwu44fUiH3NDPBq01ufxp4XsQ+saC1tL5p78Mtfj1KeV
IMgvTnuW8xPnRsEoMcrHKyvDYIDjkUHD/vM6RJYFL+bbIMGCyZE1M+Dvw00BnyX4
TYo2QjyipsJSelZ7G4alanicQKoPMRMm/Qr1IfAbtwMQuVgttkTwWbGNCs+8aIW1
zgocMsW8K7gdKafUFzxRRiDGH/CFhZUrMf9PdFaso5mxGu1UKFrFbPt5I5y1Qx6s
QbnHw2+Zq4QlTWT6/u5JSfEEzjfKuPMuQPCYQLG7SaJ7J6nD/OBDyCdIkcBRBlgV
bxb7tJ+6Oroi9AtHvJ39mrLKrfgXPY8w8fCSLfF7CTq2Zvj/nK4mkTWII2fRIzDl
7y3K2/VBmIxTw4CFNBdegvrUYU/DUqjHZI+8FeLKYCvU+u0uIdAd7D+pf/ZZktOq
rpBbemt8JxvVkLwV5PJp4kiTR2L002qvEb7hudjxeSGkdDa66nXbuB7b5qS8AOMU
pIGJkaNgUzkwialjkXBX3KOveq9dX6ZHJj77d6jlQg9u5FbjLXUSX4+UID+SDA5R
bYvzGCyMuYE74yetrtrCSuAGciq06ZiEGboS9lIXQhZMQ0tcPPSDD8H6zwS5TZhY
P7GxMnS/edAmz1E7oUUdpHHroabhXhvQ/ROMHqPLRFWkyu5+tH2e1L+stI146+aq
ufaio6QAE+hu0IQjViOWZd9mbuHdOSyw7D8yBOufh93qvC/43PmB4awoPuxhnlbD
8KuDgVu8Dn4w3SQtspcHvDEUXds0j8//1AK9ayeEHkUlXo/JiXaA7b1SWnfzLHfB
sC+yxhx37exMtPAP3iQizRl8SiY5K1vvzYTMejUrjajb6H8P5bS+cCNUCmMLGDgF
lzR71EBRVRyTFgY8+Kp8apKogCVRVEr6BV27auEhYfaBIHN5LP1pnS+xzeZPdk4Q
Ay4R9STwdjczv5UhwXBvCWNRipAz+K4Um8cnvWFvGUo0pRTJfWtT/26xUewS+95E
5PajLJBqXVKgMDq2Toj+Tl2CjCZZzxklqT8OFBuCFj4U4YSyMQZpY5kP+yOLyfGP
5bq4Ws9NWqVWSV5oc62XzSwQEa+GcKNv7c4wkv2pEh4aosP+BMcP8urNPcEj5iHr
NrFu/BnB3Hw+TEvwvkmFHMF3y3SeqFIYRetQ/wCE4N31rnclKzLYUqbEKRmjrCYQ
eM7jyv10lHZRdhKPrELhCBl2t/hJCycBd/iG+YlUbTcLOeL9Quq12RmEtvvetg/O
Utz3RNicY3BZuN4GGxeC7JxPgmIslOQdlMYmKYVxdcd51KbSeRY5k9ngJBkb3OJ/
N+t9CIgm4EXep8x3B1qMELphdctAXntVyLxHcrieYBWDBupB4YdVxP9VXZjzlx89
VED/032acH+BqNPc0KnGbeXfzazYt/Sl0J4Tg+K3Xx2u2Hrl8kD3gud5IxFduKOG
2O7mCWpl/+QHw3f96ndktlRufvyBQhangRI3aC3A5HH5qwqFt5vyHx/Or7y7jv7l
xTJ8UfoszbJCMhL5Cc7O1thr7J6oekXOwkyFsPSuIlV6kysVbLFZV4ErLdxFf/Eh
NRDVK15gWfCeHCzopUvVxskUqcNckB1Ee4K22kiEu8OfZkSsISrq4NBcCNZln8Lp
oce3ag6N5ipdxSEx6a/Pbdxxouh/sVgDoVMpxeCtnhMCCXwoZSSBzzfcXVSvqYN+
dRxFQ+IC6SMzYYM02Pq90QDPR/57pkNRGXg6zVrOc5ezT3Vdc7hZR7+13cacChNu
rQ4E6T42Vhn3xEo/BuOAL4A/Ar7YuSqDl4RuO/d9aTlWBReD+k4oofi61aqoNget
xLsj477B/kUrF1yX8ZHWkkttDUK4R6jul4/G10kC6fh5TidkKjz93JAlIiXVoBQT
2jY5+BtMZwWwWpolsR9q+tHjQOTZjeaqK2z/T/ikHF+MPps7khrtT9mQpivk/AR2
34FhglTLAeXTdRfi9W3a33vH000Np5vgRoMld4OkfdpkwJ2B1hShDHJ6wvmXvRUD
8+e2kWx6bK4wF97hwbuI/ujz1Pjvj/xuxSX4VVmMnJDgzQm0NHc24vThqX/3YGgI
DMf2GXfk3fnTZ6ul8VSzI421syIA5tj779iwHZaj4de7J9Pa1pfbkDZQYFX3C519
07Z9yRtpyOyiV7cX03eOR+1d1owICh5q6VX1fHFfiCYO3lZO3/vW+XnrG7iIVMed
8VzoGtx5GuHZv7w2KTvB796Tt0mdrTb27rbFeuX6GRWA9dfYtF1FSKREYEE2Geze
gCUdhBRi3T90PqSddXXK+oIRj2GdIOeidyu8PYhHMB+TbDdvO9xKKku3dK+Mh0fv
NlUy77tMQAaj80PsQ6FhrZmYvDoNCb9Y2ANpxh6BG6pJLixZyT7hjvSa6qEZa79q
QPxzht3dZd3au8Wd53ZZFq5Mi1jYjOqJ2PESVBDGomacnvVyQvlLgGNBnEsWa5Wt
U1DesvBUQRx64o72Yr0V85kMJmfgKPzPOZ0v1IwpcdETqecqpZoebq/AyXNH2bAO
X+qSxj7nZtpEVJeE9dCo/TpiCxovQY6dOCodzCG2Woh6yTz/pD4jCcH+wZFjhhAn
vS55z5cuRqsD+RpYqsyK+v+RnuCxNhcrQRAP52j/ArGNMS9ySZHeFKKZMbz6yLIo
e6TN6fvCMs0Z06WCNIacjUD1ZyJWypWAAUhi7vjDtAu6QXbQ2WOBXYS+9bUPxBMu
Q1xRP1ujj3VYrFBiej+vCeKCg6lWVpIycFiYwpd0LACZA7ckJ+ymuGGFXqAuD29x
iAG193jzXfVhHXfOEWLNzQcA/Nae6FBYQ0UP8o35IbxsuAYrsyHfEFSpjb/HOJZS
u9qYbIT80Rdw9WJNVZo+81fT1mzhksaYCMyLeUrO5UmNtBHiy/s2H+WoRGyn8x31
1E7XgBQPd6j6CAOjCh9iK81cS/nC6rbgjZXoSgBic9RB/OtHxWj2pfZHMreBIwex
XsQnwi6soJqZxFewjA6nNtFv18+TRncP0uDY0WgedTU99d4rvYrR7M8UjLxScmx2
bnRPNORNEd5JXby9jDVcETJgvt2wrAraoktpK1jCZ/xuI81Qh7Liu042XxMh8Dsh
p+CqDM2Ch1mvkdXRKOOi0rlM08GwGnEcw0NPTwxPwb2BJSGbuAB7ZYyxtb7sH9Aw
jDc2emP6+1CbNwOJ5mwZzh34Ldo3uTIpTkh7vvGE08YIZwExfj5t07pQ6mkeAdvR
SGJWssl2gfg2/wXPMZSk2oY//Q9E45ymRpa3Fpkr4cKtnewLEXX8+xBgCFD01cx7
25MzbLUVWgSNjsInCR/w4tkdOrh/dBMzS7j1Aclr9EDgn+CfM0zw8oNs719CRo2S
0moU/YOy3q0AXfHpbl67RREBaagCzFxLUOSXL7oV5MfGs9jn0KmLuhu1M+YCbXsT
QuWw5fWe0lz63r0rn3OEjPr4UBzzmu5lCi0nD6podDpm4i3uiChWDjD+YytlvB0C
EgWY4/kHyronwgmegZ8Gw3EHS3SdTbToaBVKVQuKoJ7srVxz8BdpfChzy0DCWsFx
56UpnbgZHetFIgHe0aZiRHmmJUtToS/9HIHZLyCRfVURTGHQ9/xXfBabII9rJk2b
TOgFBV9ofiqmFUicGKaqJiTbLmVJh9o+R0Uyk/YbSGqijnOuqe/fq1alLZnguTXN
UzGq9pQ+7/d6aCr4VKTmBu9CrWJfAeAy5aC/+WS38kKuAyvmOXtzGc7E2W7YM7ev
8DvTImhBZvuRQ11crDK6YP8Y16kGSK9A0hV28gh5cTE+k561S5C9vr66k7rJPaHC
PGeye9TdqR6N3TJbaQjEcv0PzNzdcIO0kHxmMbgDkILtcYA9wrGeWIjgQD2i3D2E
yH3F21VTWjHI/OI0pD6EDyzO39i/Pj7GJbjILYjwN0yPtI2Mw9+wOfp2nctwAAO4
iYBCz04v2dL9ryGxZTrLWuv5xDm+9ndqPtgW/K73P0QSKXKh/hncjBgCgdvZ68hC
9b/zPnu+gmdsaCCJDr7bC+9dnj29J5n3lDsiyFqoWv/mq0zsGZBOYbPH/p2NNmud
R4W8kjdFqZFu0hL1rLsbHAoWWogGRoSrp6u7eVDdlX51so75f4I6jL0bYmjbe0t6
vIfF1sX3BMq3hjI0EpBE9TAAR4Pun06niUJFXBOwvEgSb4xeAnxHdHVYozM+dFNK
KPc/JebS4KvM2GQ5GeYHyK1wGTj6Tijd1f0HtwJ+gP7kD8mFTaIKEpXHE3mruqnf
AZ7/IKX1jWwXks7AykZxiEj+iIi3Y/8D56FnPSSeY2hjL9PmVKd+X59i3lX72oP7
DN0Wuuk23791xLS35eWyifW/OcJYbev0FA7C1iWa4rlWXDxg/PfcJRdGtRKDd8bT
3oL3ag9P8RZuPVmwtdzz2fnT2GeNdQMO204OyEPFqmpFK8gQNZIweyvMK9oYqptN
C+REskOlON13Gig6TwBAoKBXD6W/nbtVF0uuphWzvM7CVcq92Yz3NoeIxALPaWjD
NIjtFfFyjOhpX1S0XRYz9728ImfEmKlUN1ZEHp8lRnGO5xcv4HJIo0iESRF4d4ro
WBuvRMO+qazKzAbGyOQWVzyEsLYO/dPUZ7VM7mKvQCuzXun7QLwzp/8NlycuDpFg
x8+my89N2tmCbQ7wYsYBoRknmEVlSbyG4T+LWDQ1GrrLAJybDJYT7Tq0W/ryNMu/
uKN51M3H3MBj5uBUWvoAxIzZED/9DclsU9iVOuLpUMRrN3XSyFbfYWmyphbWfhNh
tH+5AAgWQYaWZIgJf7oi0pj2HdULL/KwUEIcovh1IIu73wbWKZpWyt/AC3LaVLZ5
Z6dD6W7naFPpi5DrG0iNkZU/MceDOU2KoCjgUjbMzGQOtOX64DMprpB9oscnbt1z
3O/9gww7AghmgBwcYEv95DwM2wBdySfZbTFzbmZjjQt9qoStSV9mWddMTAM3cvZr
YhtKK5wabquOBbewDmkp9UJL6DpsbOfXQ+S644g/IJ2mC6AE2/CM7gF2QE6XS7S6
N5qwdatsSyQVhDvHB+ANR/5H+6tZHjGc7BJvjeUP+5BVW302BV5fCD9exPWdEX+E
7yEFcIW9qnrpn7tOqv45ndPI6VWtU/dSN44my7TJ2uxuhC1ZSoxR7moMN/6TfJk1
C/lQp0LpN4WpFevggljrgBMCVPewn+CTnpbUjzhdp62c4JciHb6jVpe1JJzdBwJe
8XSkf8/YqkF9Qb5GWrz1qv0l659LJ5AGqslgRDnq7f1nzp0o8f/RiMowjPeLN2qs
INnVONTRAnFcffZv1x+7hyLI0793k2lndHEGO7KzICt1ZNxxipazpkjuC4588YWf
Jhh0roJwgbVKLodDPSYHsl5F8eswb6Ip2rIkk+NYqr2OPlUpysnZkYSQSlPKAi2v
FWWyiZgiUa/tjAMD7jlzXjVI7QLPwmQnCfvdy+Td3baG/bp5IFbP6TJYiARPIqrS
0tOPCyXEagBkkE/7f00cstahqpKrcbJ+8n8ZOEeRyOYS0bl+2swte3jNW57P+Usb
emCY1Os2D1b3fZ38Rr/M0Iv42piQW14Uwx41qApUzG/7g7fxnS03tEoAXntHD6LF
VxK1NOsx2Rythw4jqmsYZ5Zg4BZSLhWbuC9xkPy8puduP1Dt2X5CLU1gdamQG7Qc
5qH6lKp39bM7162Mg5FwnQPoyhAQtBY1BQ70rtqfnAzbRTQEz+0rrz5u/3CCBfhm
c/17O1HD8IFoc4xn2nW30UUq1lWTLGuDuZrxPHa/pVVQ98Rcc5k7DFxNSYxM9gv7
e0dlG0OfVd5YOf6djNTqOZp01fhQX7w1iUJDmYk1WPvdEqGAKQYKwK8qH358A+FZ
m57PeLocG7miMMdkQTZ+U+9WCCtx2k4AUD7VDFFIg4YqFrxgt6haH20nmhxxbIt7
C3fQC4dy6wtTkvqlRBanHjZqa1zH71I+m54ciX80KcsKM4JwYjArlAgkkBvrvvH7
fSHMQFZZEOFhpdvhtTJN9IfKueLjb6bcJn1vMfVGfH/555mFuAiyxq2CilGr2I7/
9iGR8Lnw2/S8ovD35Iev4utlSYgJ3I3nepKvriIgigd9cwesdCUt5+/St0OSz4d/
bzPVdA7jSnLkGntWR4DKus/avDXft7iuIFenDTjKK5H8nWdLhR14V3c/JDwM6+HG
y+8WOP67gCV/Ha08VnL1sTDAViK9YNbvO+yPslosCBhuElCcpVYjZaitLcYJSrz5
gjukBVOowEgG4nzv4KfjbFt4eyN2eS7PqqfeQlr2QjWqQ0YHWy+dwXUqNglIGc0A
aq5JQcWg05xzLFtp/dLOOKfxNoksH4mXuJVK5Ool6mILUKNWMSi27cNOfg6pJ7pb
5wsu+8dl9ii9/C6/geUFlHXDfBQHEzi9iJh3/Akaf25XJCeaYlCftiH/7KSAly13
g/waxbbjYNTHuUCpA4xebnKE4zYQKRHR2O3VuPDweFnsYDbvMwypi9J5PMBDBi+v
2OsoZYHONAihkM6D16tdcRCEOCh7V7RSqlB8uEfCaXGPo/f2ydzZHCxW+A4k0y7a
4ovCAle5aqlsieeWBcEoGn2U155HAdX7uy9zt8jTvKoWxflNy6QK6DES2cdIP53z
YtBNLi8uo/LzNa/5YvMmMr9EHBVtRCrfXInUYVLv2PmLhsE5Ozef7Yac7KKSiqVd
tG7lG1CabxrPVKuOcRg7Un+mtPKFa4T9sOknoPaqtWXEinjVhlLFpqhQ0k54Lq+1
EPNc380LYgMyGMyscoai8n//LIl3901cBD+14QdQV5ErE/1R0RYSWiSegCMzHLyO
93BHTGF5HgmDFvvTAFQCD5EBBCV/JUdjVOSkOPNGnq4Aii2/FX1toJB81WbdAK1v
MYDIbB+gHr+2KMLV/zJA0/cwfisAyaxq9RFg18J3u4EmGvmtp2bQVj8TK6b7KK4N
2zyFwE7uzyXRjiEtsMsFnlwXFDo5YWIhCmhZDEQ5v6Iszdw9FWY0SK65+Q+zhWw7
5wf8V5TTt5C4xLcNWKIjLt7RbLyKodnReXNAjkc1k9xhpk1Z3ZVg0Vj0R0BRYZ6Y
EuRHABbEH0v7pjiOQchuuh7iCwvANlkvVMPR3+alGNXY0UmBCRm41fhyO7VoVX+/
RkusNh3dpOrC0B/flt2l2ZLslNMyHsn+4EGyT/dI5uhCc5ftpLzG8g91H8qHiePp
nzhj/o3oPtY7Wqng7sYBc7O9N0CZBE7M4QKzcsUcqqDAQZ0adBs7MRyhRLtflh4w
Pt/AhBDCxWPOKUSuHP1xQzq/mF8RzoVw23aU8qe705uzXQbbb+4/Hu8JpUXkyL1v
KgNwt8eVl5KezgNx31gWHv5ZJjNhg6vgakb+SwM6fdVZ8UBg7lym9eaOM1Poc7wO
bLGyt6yZ7H2YIEBHwDCgaIqXT3czhoEhzM6fG4brdpX5mHiWcFWHcznMmxrjejuI
M+VOkflLfIicxBQR5qQk/JuPgnNqtvZfoC8TwupGhuM9FC7+MespQNLDR1V8VGjv
eP1ju3rYJdHfk6uDXtEdBOaDoUE+v2RP5nmq4nX2LCAH10FVUTpOogs+FzYtP/QN
vG/8Yo49Z2GexokpZgXHQVdazoS2e7tqWiHNi28dervGEH0+Lgaby59Lom/wDpSO
L84fzzaEWlZsKYuVSCSgfyk8TAxptzyNtoUcGFPXQj6S1VXA1CDmkIuDevLM+5h/
NUD9cMud/qwSCiY6sPB1bu5dNmDAKGrWqVaaadI4/Cur3n3xrwr3w+Tjr5vbgMcs
fmXMcIdLLzAizDLS07ZIZGmj78ifyaGspp+8HgTHCPfQ4Hrm+DbpO7zkoJSWg8Re
g1PM4AVQwYAaPBBwYcch4cyJAfkD3uD1kIT+ZmeUy1CEvhjr1OMNcKY3kOzvAlDZ
mECw7Hf+5Uyad5IJ4RPu0+NXGomoMyPWWyMCTaoHfstkEwX8eSoy4hMuKH25cnyo
/WQovMbPbI7S46lwMSJAYE8WQGbSjFxMlnaoN9X9fvHTbWrqt9BVY23oslGkVXfh
Zm1ctMyG/I27jrLmdZuLH11uV+r5RSMs+lP2OEQK49VrNO6oJ0ZipUvbg2N2chIv
QlhufZ98CeZ5FXVejfNHfbwWUZUV46rDkFiZadruH0B4i+oDlxR/duhiDcSIORTh
YA6e/t2/N8me13a+AQ8ENNWPJT0RThvq2lcSHD9iXaiH/Ua9M+3xuI193DXELCzA
XhCWNCvEHe5bdaUzFv065mCV45xsDNSA+RXfGzWsZaAx+xJ01bwbsOpCC9sSGSN2
iLEoL02JuQxJ49Iyf0LiVFl1E2m5q9sOmzsy/DP7yepf2EsbKIsbb0WhVWbE9cbN
CiirJAH2oaknAnUO+KjBGMYFz9mmUnYPGRpzgNYKcmkEmplt01zvq+secDQ5ksHt
QjyJtpijo/rOxufGuZQKs0PAfoAzau0sIhVbJPnNBD/JIJV/06jWhPcCGgJkDEis
UnpqQZYaXsZdNu08tpJ6HAkUnq6Nt8XLdjI4ccTwp1wU6IhVt+4DWT0gfV5WTaR2
7aOt1E6OVn30ICRu3AxvBi/0YVSOw1Fh8GnxWHbU2CGv6BRMXfKyaD9odsA6YVhW
hlHbWUlsRLPnkyzGGAuKWUGHfprq3xjFeD3Z/V7HtmSyIorpyxqNHiLkB7TsFFiI
vye1tADK+LZnwd3YnLNWJ/xxWsYW55W1mbusE8PHX/LUrW1PWZeLK5t51hmsxHhQ
3w9ITHWEJ0vvlHWViOfVYvMltnKoqZEQY+uosj6q00EI5rdwP4dql/O2w7OFK6P5
EKH+cGuetp4AG/7XN5tV+Y6UfTn9PwEuK7KeFgTZJU18p9R2/Dby0sSPA7q1QqsH
1jH54i/EJZRJAE20Tp3r6k1aYbnKmpckFONa461BqVbv4l2bZznOCtjN9Fie/cza
WkJkEKJu1cB7FhjlQhZU0hajcSjtraKdDTfHXJz6uDBmcJjjMblAdsLY694/4nDX
axr4DNzM8E8E1LLCwK1SJL4SHPZyzriTwObvJQrcG4zZlMaJM01FeV805wd7E6UL
s+H5QUO1dKnWFFQoKGSERzd0ryLsHpq/LvYmDfwGNE4CJ5WcXlkn7VfAaVD4YK2K
ywm8MD2GKB81xS/kq7v8zAbF/Mshg6fatYBp+PoP2a1EJ8+4no4k0WyYrXqzyGA6
GDjaYNa7/ZvH6WUjZHPYqnzQVj2K7CKwfZnVOCVkYqMsZEY7ZIhVec9x2LFvxgPo
2u4YqvW0LlBHoTwyd6UU+ukYKM9drMVlNtnjEdsCcZAyDcAbj8AnjcPDnTXaQgvs
f9NWnhh+MqCO5XWxMerh93cXo+ft2AR7pcgECDSDjQ7VAOEXvR04cnBDMQTrhtRO
SVsiH6uXthbdrXJe8ICmzyZz0mJix8xL/HW1zotzCldQOP+DHnEGIe1naFT/Fn9d
pYr7C9lVFrcZ3Njlhg4aohxOOhd9EYA6Fh+QiWunPaPdSw9u2v2SyMhkaY8Oytxk
D1oHxcrkuT8BxRQySimYyjkRxHQ/hNvP3U8QKEt3j36de4p51FVE92mBdMIMxNPN
g+mILyTSeuIgOx8YslspuX3TnyH/WGVT3Rav0hFoSkCUnOTOK1ciM4ABFLN7CbAG
er/UzyvMnx309CiD3gAupCWX0TjVvaUyX5x2f9Tdu1fhxfESYUf3a3uaIoTrZPii
uruyVoomZKaOoTsvT2SrXKEeT49xRQDZWByxnO3mFUR5AMOFEbxYWD7+s1gZ6p39
rSlZhq5JP3kc6Tdk4svyIB0YOLF4nhuvx3bOXdjS6mcB7CB0Ac0IjqG1oN9lamF9
9UcDEDACYR0bxCx6JiZxk7DJkAFSAh9mNag6VKcVT9fI5AESoaLX7wYwGowPwnPG
TbiWWfoeizNtxOn4CzB0D8fwnfCNDOb1WM6m4GR0BNqiiyeRx6Fppm2lyQ7V4wWS
MePL9b0qG0nY5XXoBp1TMV0B51oYTFkarDyD8l4733fXiLMOhyTu1lhA1Vxiqsbh
8m+07rtYQw3qwuTPaYopl9Ia0h6Sb+LqvCkcHtO8+nJjiMHa8579JLLfc6vIXZ0I
rzRZ+vB+kz3+4hfl1IXSEBTvKMKg3e9mSprGyC6VHXn6Q9/NM3YthC8lHaXV7sDd
hx5fvv6TsAjlDBXJ8skoJIkBYBxZZO89l6TjQMh4mKj/x9WVozdmdo7QbTqKcmgQ
j+0I8cYebHLMotbbnU/NymUx+EcaXi6xGf+3/fuOxUrC0Q4R6E7VXvxR+6bmP5k0
ry4ZK2235/+leoJywJHp9DlSan/Egy9xlsqkVzuzzwWxDtaSnLS1qZtNJunF7+si
GTKy3xbxaZP0o9s1r60TjCLqd1DjUOT4dzSm8M/6zQ9c+wPT1ES+Qy4NOEHLN4Z5
wjrCACRGe5NFsfH3wKsa/CVp7dgevY8KqKe4+ZCIjMblTXwPRm8/c7DkEOamC9zG
0wv8wINZPahWB/QdLBzS1RXRkzHBD/FlzSqLT6t3zdgbvjKspXUETen5vza6kdN6
G5LFLr6yCLpt6pNc/Was+Q2a5dwI96PHjaD/P8b9LkNxe/2b/d0C0C45mTH4RyKB
h95M3Aa8HhOOyQJajtSCvGxDIq00k4pFXt5ZA8wCH8HcO9+qXzwH+WuaNWEmUZya
ksoR6s7mdz9z6mbvjPGE4ZZ8OAb1pR9rmrhbA/tlKrsBWjqL7eYT7Xn9LbxKN3uX
zlGGJ97rZ6A+x7IBwYFk8ec89qGLbZhu5HNI9arhloD5k/Pnnby7bPCv5vnEIuiT
Fmpm08xG2PfuU8XIIsThlccWn/VcnEI5UPB6U00kERd3O2U9eLmB54ZppDgPjnnO
s2HZMdSo1sB+1JxUW2XjlM3s1dxbIbvTja2I2Z3So77TgCgvHa3R41sDE+2ZHU/Q
HyksriEjrAa6pymaNQuvAZRUjAjo3A+aGCtmbu5XYmkG8CJnEns/oDrcYjEMwz9f
d/WUeOJGc3Umf9ydopATH9EXhNwcIblzMtEwOaVUlmrAO6231w1vqomlitE0Z++Q
LG9SonTUXZH6+64aixZsOOjOPwaDwthIA4FP+KOQ/MPY3M0zcremDZKhjG+AYFLl
5/MYRaeLcixb15tr0eZ+UNlMVyt8lP/ouoLGmASyHxWfw2FQdWrTGKgk2xlFhucq
VafZZ+gBnL25ShwZZo0HAJ2Ikbha6z5n8ejwe8MKIjsU0UFij5SwZT7FoSd/Saca
AXoJbY13qfaC5q4CvagcEvAStmv0Hue9Jz6rRKGJz1i1VisE997cvZ2dXITVclX0
JZOTF1KBOtEMDjsxVvDtqzFGR5/zgN1CHydrT5W16Qm940UVNE4NfUWx2uuIh3vx
ZOmaWQhIAR0wsB7kKLM6rbwpXutd0s2maoj9pxj14ZIrYkgVQ4Itxb2xqi2yazmt
FNTQCpj4m2ZT980M/COR6jBS/v7OaKUiYzFOJYh4zdTa0LXyPuT9hrGM00EBwQ7g
+wicqIIrcRJYniiUyJ53kOqvh+bAacTq5OWbCjuFIxUKwAOAI4J8+ecTVWQfYvgM
IYPelr8nPz3n6xVGX0wYsQfg8ZlsYO6J0rD8l+4NLgfoZjmbEbut+TN0oCGDaaKM
4n5sU0ZlR9FO5oaDXs8jEdi4ETRAHSqMv8x1o41Zfr0z5RlNRNKPO502UzOutAl5
aSL2YmaG5hgNosTXVN+CKi/UfctNSz5Yte1Ss3NuD4Wcz8PoAvmMv6syS4DWNeyn
0BvebSoaR7Wov0zCqar+HHsbvDc7wCHdmZ68vMUZ3UX6FmZ6kZkkjzOwU8UodDtV
OYzkdkbdaL/zGW30+C8FpwPyr0LQi50fKUnyGmmy4iMXF6SCWDSxhMaURAMO8XcB
2F/j6YqAk99ag9F6GIxdQWpQCahzjtgAnDFSJA5chnmxZt017+aoGbNa6qU7dK7s
901w9wg4S1m1eJMV8LP291/2GYTT+ct8NtD0etB1ofgTJSa62IuHTpJuXsrnIzyh
gI1XGUtilGVnc+d8bC8yP3KoWlUmN4R7eb54Hl31WgasKPkjhOVbgMOvoraTCQ6I
sNEsgP5Zgoy7zng71Uw9YmBoGRWC7cbUUlxHNwHl/Qv5GeAtwJSsI19v/UO2v5e/
VdFp9RF8IVYkYQm/gMGW5IM4hOXgsovFgWGlVpt8mAhmIaal/JyjtqyvDz9ZlIaa
LXGxWBy8xoj7Q82mz+9G3ks9r/uZpQe1A08ljZnW1rf4NdQAHfIh8S8+9cj1EwPl
fQ8CvqGR0FrOkphVPER5yVgev/hhGbzlMG1RD17fT3qpfRDMxDmjNI5pzfKmXIf/
LFDUVZ2K4Tqhzn//Wmp1jK7iTWamAzb1Kk1d65j/1YUwj4///bhQzb+bQ5CX+95b
qDXQdDCxARzYsWAmsfc1nkMMPY/1O4DzvbhcV47TwpnzDXnlOF9iiGohoelgl9hn
9+A+j2IfOS7s5qFYtIGT417n9468ulmoewqESR5HAFIskAapTdBSEzmCbjg/MaPU
vUSMOhQ7Xht++A+7lEhHdGp36W6r+Ewkg7X3D8OMpJZSCMtmQ2J3h01i1OR/ihhx
EkoHnTxR1r2hACQrMErpQ7vyvyoiBvqK81oizYkkK+7TINxaT7cpBCoNp6sk3uKP
fanFPDXGI06WYJ2hUCHKdFq/xdc+/BjpaG+vQ5Xbv/FL7ciwvTidHzIhBjfORwDr
8+O7SC1dxXldt0Ngx6qFci5DUeQXzEa177Z6o/oFXDL0ps9GglWZxso/1jtBPRoS
ziba4xZ/JyemolQb+9e5nJBYwamxHBuykKip+8/IGP7+U8XhNIeqUFw50gCkv1HU
9BvOjKiLxf6P8IcbFh5MuUFEY6h8dcHyg0QV5/AFKse9CocNVeUdmAEsnXIsBZNJ
PUdSJgdwco+OdEuuY86rzahRM7PLjlOomvzvEwCU/xNwbyXTry8n2IMv0e31q0vQ
vyBsr6qKnroPlN8EDSct59O46mLt/H1tPtPtWb/DmyGQlsgUpXOT8IbtesT+yzkK
OCbEOMOwpU1tV/mYXIW4rFD2+Hqt75GV7B4RwzfcZ5vr0rOLBmDTv7canF5mNfpH
up7XhhH32JFRDPAVTCNzWjsCTup5P9eEcirgGSjTEzRVV36gWZyKDonEvSKRAHok
dmCPRipLDlZ9hwInViQkYF01hL4znq4KnqHIUzScHaykDlqc/S50J91MKjQ9eSzU
Z4hqVo8+1ijJhM8JDLV283/DkSlSAWkbNeg4aunjQHTyoniOlD03hDAzdpPmuj9t
eVO8Y7wPJXTpKue2zZJYfAkXUK47DeIIFHOmdB7v3D8RoAiOQS/rWjduByP56Gq4
J0PA1dorFq7X+ic3ZHf9Kl7iWsrXM2fAyWAIL65fR+J+t5B0/SxCwZUp24YFLnaq
TaLxtwjycteLVQy4pMxjw9Nk3om3o6S2v25fqDUSv/j0zO7NQ82lhB0hFPE6TDEn
ugR5Dm41HNuxgJMB6p+6wrF0TSUGMDEGmoCt1gStISTO+BG/y1+MbPwOs+8bppiN
YF3SJ2yCQeaDjCb7LqZPpCCECaL9xY83C+WKXW57X68dHJ7iVQYDwJN+F+IE41j3
N9mTDfz7RPNPRYr+rA0MJQLcBgWaUcPX843/8IX5k7CaH/aCq5xtjPByHZMdKuD9
BEErFcuUo8sTiEL/ov8Uc+VnyMsyHYScFlfdWLN62LBCGq6FG0bLTPcrqZ9n78mo
YiYtBIjv1NFB1C7erbOULz5M5mWzG5StGdlYeU7bWz4egmVgjIrfvZslg8EzUDK/
eUzeh/nkeRQaKKRBUkNWGPuomfKXTTxQUoVzRClSje+SrOD7zY9P2ne6T20yJNq6
L9mJS4jpNmhTotk7ubVLw8vq46hTUPGvBnRouFFBRYkJXf/amsKRGzv82HEcJ67g
urboIJO/JNa9RuMGft+4+gPqHAxXunrZdts5gJdvi4KDrP+rb9Td5VVU9Tk+poWy
GHr9gXs8UF7XVSM2Fczs7Mhu6RtT6wi1gmS3dRSLQuWZL1Q1N91Qio6N06Fs9bWi
tmz/ZYvWUq0/E8N3XLuhpjiu6ImEUI1/R15geUvgzR6wWRgez45O+DzqzC3eEOxp
DQQEYSCEmhejRbpXNSpnSWZ5YWnucncy6LGe4FfrBaG0+FsDwRax/777duEL/MQX
hAod3pAhZ30uxY4fwtgXT9guo5eP7BrvERHmC20j1F5HeJUPP94cGrSiih3FMy2I
7PrbonN3iAti7JHByFlu+rfBiSimnlTl/c/NQDhBc6z4LWHER81KRZzt7li5IF1Q
NGd+A+i52zqSMGFzOZDVHxkGQMMLvT6rbs8DVgmvIlzFXCeo+GTvt3Y9bRBoQayq
v9Rn7xVRKnCj5BmvxDZXGt+GQaWnXBCG/iyXk6z7l9XP9CRGlnHYphglocuuuzbX
I/1FS/wA5hxk2GW3YCtuRAInvvz9xGQ0bTk4Iep9jdIuPop6BqHGw5xTZ7PDEd8v
NH8wJ5Hm32PttAcatdrF4FhxATjZpiMG/pQSzkwBi/nJMo1J2vXPqhbyqmGR1iFr
SCvScvxB+A5jEUh2sesd9fTR2oQ3OzO+KHf+1AyfHFZojpL8SPTIgLw+7A3ETp0j
g+akrKfeH2gbmmLF9K/nWR5VE7Z7vHMOfSlrk3Gw+yS8IUoepP411WqUhrl2LpVY
viWRmSVUjdlQ/zFZOxMD8xyR7vhlVjueuLn5iEVmeA8XT8FZ5ZzrrmXU0NIjgzmH
IEGyZfc8qvYDvNwZpVilk0K/lhjFcPHhDC+iX0uY1x4QQeVeLqZwTZ/V31XWgtVR
EVIhWpzb35/6pP8nZoFPBCvyZIKg97DxYRgzdlBaRNpNR5n7EQ7LasPGwFplXakP
DF5xnQN7Ltbe+OLD6A+3aLgdtZG99bOR7JO6BzQfuatHm7WzoLDWUTJYUhnhuXH9
gQEVS5KxL+fFG7qnm0tTyuCDK3NZDJepbaENvfNWdf3x1/3RqaFkRUKhLxooa+TE
nXFqPdSmfxl7kF2+nxMqQS40Y/RcIdaqzlgGLLrW0MnnCghYR58Exmsr14Kqmi1I
6QLaz+WQda9sRcyXxagQxOqAnv+zKg/prg6YDMX1m/QFmev2sc5LDAnOebfUZzF+
OVpUdp55uGV4ZLX2HpCXeMlVnGH1lL3Z11Ijkhm5R6INlvPzzvcWqebw/VjaIQDD
8gZar/OhYynC9yV+Nl9ciCK3tMK/wFvxgqBiNy828ssbTraJIbzuS/eqZh42Vcgy
W6M9veRPN1ERCNEepmvbH/Yea/ZjzKz5ANXoGZWHtQNICPYBUc2QMcjOCHywhxMx
Z83CRVxqAIXamPIZXg0CheyIAVaPvqY2T/LoDOSiOUYnDzt8LlNwOxModlnnv/qW
8gNxtV3GC9yGf0BPyYRrWHuJiZ2S5Xn4XsqQbJb4Icfx1DV/nmWl+oNwYdRKPu+p
dZCxP343jkfpe1SQESI1PSkOBApxCBjfZX4ortap3kRJOqY3n9pYxk32L7PPUN82
nA2a7qAIbMuYYrbyDucabm5SvfO5u0Bhgf3Sk5f0sf6JKaoIYCntXYLaE/AjBOsg
IV7JoU6XgxQuEPaIuxz2Z54Ih8XXbqBIdNBcRuumw9jTRT4ak1GQJsvPe46whLMR
3nmrZSvRLcnkANGDdTRWoklHqDr4nwwwbqkktfFIsdoZhA05/ygfgUXHwhtaxVYV
iWWXeTVPI6bOL/kx8cVaVjCAYbfBxWeYoldpQaNBxsP5vvHSlKtoI68uQ49Vn06P
SYazNEGcV30ncHTdFJRI22JwFitIlbSVpTeB1+K237Y4n+40P1EE3sW8eIh9QKZK
CpXkKHWjw1mjybHUJbdymVpZp8aWbZ4LOblQ9R+e07DL2CedSjl6+VR9kTbelGkf
v4zHA2PJMqJlCEFdTOsXBkLgQa4WOMfwsZbOLbC/V3wcgkuZuVMJDgFRlxybMtG6
2XG4jr+7BZlImeeZ41eQqDCL4mlCLSyoKRX5p0zDBi1qImciWdYCq1Wm4AC6Tydj
tPSunDxqlRCxq0vOQv4gk6zW+Xqw3zrJYu2wRBnsNTgEtuaVdR4AT3z2EmVqhP9B
vDsoDAzc6j19IbxQFQnJEaRO2JTYYkCtH02/+mh71jyRUB6S61g/6Ky86ykku+9l
nV91BYaL4Aojx5JPJ/mbJrop6Flf9bXUT3UY40nG99IS+q/tjjSUGNevqlQvriOa
vZAKNvbc+FHZsv9QenYYxmwKpPxEkcbo24N3inch/hjISKjmpVihiKhtLqrSovmC
UYX5SxwvXJ5TakWepRbyBRaITwj56H/P1bzG+bCaMAG0Lfk26RAKADcIe6Q+RSOB
DGT+AlM9CuopGtzZAKOxGEPdIz36VVoq3VePwuNm94ReOq37ofLb4h/MOiY9KS7c
AgDQPkpBpKQlHTWTI3TfO68j0HB07AB02ANtvWPZvzEk2zPChlQDpFL3u+gSQwHp
aU59UfcbjWoz3fGZrLFLRwpMe5FyXStOVJzR0bcN7Y6Isl3a/p/T3SmMRuupqeW7
dheOkG5eqJAq+jsUZugZekJttIf+0+jqt8Wmn3l1Kw6rF8gur8k7Sdr+e63qM5+f
8YPxZsirvUizQn4sScwUXb4ZL5lZ0byYHIB4RJjf0K2QaYjzFKtZFFoalVyfv8Ld
xZ9z1jHWz/McGXghfMrTPdGtbKNTn6D64A1MkNXT9i1V5lmqgSjLMdUoNqLq++sD
nSAyHGPOVlWLk85JDUXJ/UARAWwmMOaQfBSg55LlCSzA0/s5SYHkDDgvwN1gHRxM
9W0Obau6CsGO1XI+OsE/LaohA9SOae45vSXd3NPKiwmf2L24GfHylSbId4MP1RXr
eT6hL48hQsPLKqizzSkgqVZDvD1s8HEgCrLI/F5EDMJ/z/V1ooWlSuaRI9ytK/w9
H+pYp7n3wG4tNE8fdBeSgBCe7okMJHS6oAo1TV9asYhngLUjRbUNj1kXG4/0iwJW
iW1zdeLWiTZawoRhec9nA0igZO71qgIvHuiOOrUIOUkpboCMPlWZ8Ut9jJ0RkUdR
Xo2IXdDDYhWR2+fgWGZvS/UrX+fmt5WIcZP5T0wXeFlYSmoGVI3C1kx5uIeShM8Y
JEUVbln4TM9jdPuAuskKKm6ije7qCT4bFzjn7U16Hdf61KmIJRwUZpjBMIcLN9by
T9iDVzkbI8YcimrUyBUxSaDqJfQo6r33Zn+oGctGY48zA6JJamDB5JxmrPG+wYo1
VCh7EcOYpv1TFNxp4jdezWLZYpjd7Rr4Zg4l0NV3PGIteaVWE/elEMRWKHhCRxJ3
T+K1XVnVG+fe+GpaVnsDEWCGBYH5p5aC0wclunPG9S9bdKRO9M9Uz6kfZb9Sj8tc
ZLKGoGXwLRgEF45Uu4gUaGj9CgKKh3JzEF/g8LLXGScHfwuoHLiEEJcxnIhXwbGl
+WkCrR/J5bOAGFDkWTklJQ2xovtLd5jEi4eb6LmtCKlwXUGg8/gxWAm6kl4KUtgw
VzR/qRqCxSMZ8hgmp2NoYOnaproT9eMyc52lgi+7m2lRwFyg3b42Q4Nrp8lgH00y
+Xi+9CNG89Mra+7dG61br7Ovn0VVQGBvlkNoYARXMwvy791MloKKidKeo64Gxp3F
t32D0tjRj5Hl51Vuj+QJGzUKf+suFp2T4bQsaHSkb51EcX7L0GLaq7T2Jb0sfPD8
lHmNEJoFYR8joUMkLzf4SYAp7E4zz3S2J8dzCyYEQlAzL69bDtXLq6smKZU8ebff
MDqOB9x7a6aA/T/YzQpl98GlZU/dF75E4DesHXNeq7qdAw+C6FLyB6PC1Cj46m9s
GLxBDIvF4Z7FySnbjp8mUpb5IqFR18+5SKprqft/gLLIW+csorswIw+oDE7hw6Nv
kSld7aDVuneUkTY6LMl/th8EseN86C9OGp0+/GHvPJ0VM7SDDocNZIMKogSLRI1J
r3NedXSD0B4CyEjphRzJP4DKlmDy4z8ryCvLyo56cly1W7iufWhF4UelDz0/auP4
3GuJdo/LrbHDUuMEffK1YkuPSBOABOWSwR/KeuRq4ea86h8OMgdN5qnpiSajGw0j
gkFdVrHiCc7IR733FlAsdb5vX1fbPny4k/WjtF3kkBn7B/EsD7mEWVhQul377uQx
4z58Tx6PFtVlJAsiHGYEvY9gUE0XfUUD+42FPFAai6o5SySPmk/x6guiya9ISGw+
Pfw/onpMOX4ZjACoOsL6lRfR9MZxY6P1uWAo6dr6SAg1MXLTd/d3mTO/r/2EOssI
r7fZqIVCW+YWZsQIdmrULIB3cWAaK2826REw+gKjycFxulCDl/e9EmHw9ktwlHS5
0SEwTo+uUsRfBcklBakXfj6cMrUume78KBaavGQOTZaoMTWqeqqWrU+XxvYgq10o
W/nXIgVdYDZtwDH7IRD8oVKTZnz25BxK/8MXgA+ZgT2V+j4ci/sGDCoRTN6cLlpR
FasYAeW6xn/CeUWLhFLDyOzYRRvTvMt++/cGHjI3sqd3wMc771iwJMnDqUJzntiE
o9eYB2oyAz7/8nySjkLpwTiT2G4I3r4hAYF48MH0kor+NNN2CSA2aaCtOMr+iO12
PSIQZwkHjWtfFD0FSHsU/PcCXK573wBUU2Whu5+xIBGcggV7MQwfvKsVusYdsc71
uiJRzxchBbIK600nLojm5dyWXw3iowTkYr1Tj2NwBqC+B1vaXn+K5KZSTYhR7PpO
4LPPzzfrjTLht3PuKo1LmAtSmkTZAF0wXWBz8qbx0GMWUAcggBFtEw98o0eYu09S
AJKUGK2PBg5VXRSZ5CUBl1FHHCVtac3mcY23PpI8H2KUnlxFl6X4FSlXUpT/qyar
ee8oDjwkUfPQbNx/Fi+H/YbnxpjgbfYcIm9gXlDkjboOea1Q52lPTx2lHhsYu9Fq
mjszJCJOoVluKhdX7FDQEyWUhjwgm1AlXxSmgX9/bpdbC+NuPx7eInFNPEnvgJBb
Y0nqi1GaJq06YUit9TSSdENg3eE8YlE0vqlq+z/qQDBbtEEltYm2AnM+F5bdNiU9
OXQVQNRp6p0rhOnVMqTN/M0KVzk6tSsMmvEm68GYOQxbG2zZCBYQnyf8UIoQg7o7
DAIiQAgomaOqHDGCILKauP5vjehG80PCDLOs7J1XK89CmEOzNW6+VLeINcJdaukc
oktSb5bu9tTbfvckuvNUMmRdXSh1MgyzHfKUajEAI3UX/E5LZkiiat3eRc18FjUL
XR1P8ZqPYs4dKQksyIP4aWHg4sw4OdF/1leNzzapUgiXtlF7dDbvmIOYEYIGGegR
IjBlgHcO7HYkLn3M6mp6HkIMiRRh+zN5vjSTImH0GLmdhckvxdL2VEKOi+TmMx8I
K2nmWWeKIGCmKCTThM89+o4Rpg7oJZotF5bs/C8lNpp+LDQgvN/i3aI0V/Ufucck
h6mVfV/zs4zvVmNUCkzVS7xjASuU+zejFyQElTrtc+JfxOe4fqaU/3udunJq2ybc
2GMyB2V3ijBDkPX0t9UdJHgXy4QFoSkjRDDET+20Z4pH99ITmrUuSjx67V300Ib7
Shqvv26Du0DdRYRhq6ftw1Z8NQJ1TJMRF/5RTDc5qt0ZwFmZZs2ItrA504fK4ZAc
DkSZmoogtQDgqY+8qGrZNK1S7ihrIYPpRbkmZND97G6pW1hq7o3KQmXmX6shY3Ui
+MFpolDO2EzmGGvk5K/7L32Wx2IxuTnduuxmGgwgWicZimt9qoITpAtkdpPEaV6Q
ovMNeuIlmPqDoJuXzMvswuvu/bmGXuOYY5CGkn+JxQW/XUv8sO8xWWPHLqsHiBQS
ZeOhEleLWYEec1Xk1KArvifvET1MROArjtsAWDZAUuee4Wcf687KAu23TTyN4Amx
OLJZRSgfykjDFQF98jCXWZS+aTEr8jMWjuZGqJ9h67GBD6qfnKImrFgGkod9H2D1
mSqmXNSE1YS65QR6gCWDhPBHpe68JsODQshKj8QXRSYHOKRCVOgfBLwsIe23ZkxE
uxZ+kjpFTD5ME5PRTKsJfFvO53b0Mc0awqfI+5z4u2NtkQsIXRXiURHT4G8UVjHv
Pbg0Oq5ST+HmabVmZOK1EDeeih2tseIo3eCF67lwXeexQ887hkFN1tJL5a3AEk4q
f8Bac7EY75lttXsl7ez9Rae5qMbvGaIsCr6AQP48hVTqTCBVdGuoHHeuEQAbhARH
X9DZzXqO8qQtQQBs1HMDa7M/ju8G3y/oMiOgYzIsMTyacmoSEnBa/KsjUNAuuDOj
x6c+s1fZH6kpUJ8mmfmNiebCKSYYQmVicQevVbLz6IXzTmT8ZN+MX9tp3+48c7V9
mspovvjscL9GGJv7f4xKY52KHZgPxUCbyM/BBZru7reL5vxMN2e3VUfTpysWz+tr
cKz11fplFqmZHw/4cnTwj5nOoJqFWyNH3epzzMm3r8mpcJ9umpgTGVkxaI7wSd0j
tkQIoQPeWB8RBgpKPTihPrN3i1lJ493LkNuUZQOcALCsZJ+Kzd20qgJQZJqkIBve
jRokQYEnRgGbRrqBjxIVP+Lt/UwZf1/hmmQ7VYSkKEEpJb1RlweSMvqHYt9cQhos
LIdv0Ychki42yGWLstLGfuV+RfX08ohRlscloR+9ziZBnV4UCZ6e+EoaMZZSCbYY
rXlQcVi7OgtQyNTr48qU73G7mOP3P3SAjDklps90Q8Klq1CuNw6wVBEEtBY7/Do7
H2UGRhtma7Vk5Fksr0F1t6zXQ7EIUxSDkcSjUVEYJIHp3UXZzqHGldNskE3CG2Yj
IUKwdZe4NYCRpguF2n5MtSFZAaUtW3sUJ5XuEDuotKgGJlmEJWydjOeqQW6SHWaW
aST6J1lAtBCjItMD6JwsyQAmUlEHqhqkrzp24i13GXGu+6lgq3oGzpYd8XLvjGSL
8o6cyMsl24kijbNebUC6arM+AT2DANPH2yLPCkRFPFnh7kyudNd9+LWsjzo5mDs0
9IlrOih4y2Z5odSC/PZdC8hZECqKuJqMcMn2N/6Oy1P7r6GBz9lyVXUUXrywKQ9Y
42epQcRw0Si1YBJm0J6tt2SN1wCgYgkFIqSv9MuNNztbQdTZc6a6WNUXxyScvGTu
h3UdJbofdJYq8r8Wr/fcdIvFhemDPm1qz6MwauZ17DJOQRsENdJhKqIGq3cDsgC5
bBR3/u6h6ZjhmbqhvJuqLeeLzn70k7PqFC3+AjDJfvREubTmKnF0hOHa90GzB+op
iGGSRdeMdiqFYehLL340H8qaF1bxcV9y/H/zFxSH4LHx7x/e9LEiEoLHKwikz3/f
+P6dcbczkK0rfE8IKKp8scsreux1PUGU8CGLJdz1fNwKheHlfp+RCgBM/x+/ZIae
J+fYcBaMsFLA+9V10BToRg8h9vy0BEn48xvQva9iYOWRLPVltpeJB8cob0LVxRGY
05xIF2yHhV4o43lo5/GGqeWOY8ZAfj51bcAS0KFZNAl85AjIWS1yrJ/E42yzMlsv
DKIGXNAo9OIba9PfOuM/By7plLtSxpzLXglZLF60S+5WA6KtV7InHGDKCqeel2eh
qHi0EnBACwK/9vNWfB7PctOVsiPOU+NJ059gWtWd8fZ6j/huc83quraVdiAcMW3W
1IYEZoAgCpc7TKINGO9p06udKu0eGLqxAYnPkSJ2nn97GEuxwGtOf8YaqJn00Wur
8xDrb17m1K8SOa+xlJWAQySEWF8GO1ijo7sskVrzIM7n1m+3CUzbEi4jTPWb2Se7
5cof8OIl9O/p9aUnDTvPX6AjUe3M3vxpfjswcUXhDElZS2ClF+L9zTs3bhyVnrAC
Rl9du+9UkP2HfSljVuIwO12KBxtghZzNTYy9XpwdrEV6XAiXRbQfVP9MH+T2qSg6
wdZgTEpjwGlgTcKlW2Jobs/f67OPSDpMltGIBu1kcyygIjFkd53AdiwUwSC3Bwv3
IeI7KMrYG+7NDMaowTO9KK83tQu8b5prKRpXz8RvEf+39gp7vQ17PrFb2E8EH68K
kIaV78JDt/qth6Klelq/qHhNAmpjr8yQ6RebJeU2xqS4DBdja8KbvH0NLsZB1/tJ
7vny53Pj/6aZHEkt52JGOYDb4CBO/Ei3VCFlvkQ2kydfSmJah0Dfb5ykehVZwXHx
xalIm+HDo2NToJeOSsBuw/sSLzGtG5RGmZfSj0Em1rK/0KL7pnZVWaPCFBxp29xT
Klwpy/n6Z8/0yNtzjF+Gxw==
`pragma protect end_protected
