// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:19 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ty+FrHQO9s+wNxpiAgkCkiWhyhqB85tYDWgtz/HfLjK97pxKbFlOG9lPIIJpADHi
XsQ89C0w3aqJk+CQvsCPq0Cw7oFrN5IGBZuiGu9PE/QhB013juoTJzxTcYCTgWAI
WhwRPG4Ft6K9RDDBYvGkg6//Nis2/JmtqqzwSGkPtAU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13584)
naWKPAnHcZVf8eBD9/X6loYhpF5sgdqGzRAeZI7F4CKr7ZD30QoPHMOLywXtHd8l
Gx53VXQQfT+LonmBPLG9unt1jLXyABIe9IXl5qGxMPcsghHrwQUuyizUK96xQYz0
fcmDCzwVq0WgK0gQHG9tAT2BsQKau+rc+2M1rcabXc9xV6B2A3e4J+MjwMy+aXUd
B3W1TGAlXP97zjVQCTIbdPxCN0+dkQN1C0zNPzvbtHJHUBGcTLZF/MjqXDbyTB0Y
BSoeXy/0b/9O/qR0kP3MbcVcdl5hmTqBu1H9C2Qk/NV8S7ZT9mzavW340UHx5EZW
CDy1ugwGpxt+2j/3I9lNv1+s26GqzjH/IpTbJHqwzXKq1dNvTr6RarIDlElyyJjl
kU1RMXv1n9pzM/CpAG7yFMurutDmwj/WCB4+BqHKN1AEFlR6D2mxZBdT71tvFF21
9FEKRvQzl0NIo3wqTLSiQqUBED/AgrgU3bXAyye6g4iXD7ksY1aYJZ99zBJHFKUq
/q49X2PrnLJ5F+TwvJCG+z/iPu+sYdybB6osKkl9oJY68v1jzybFRBMk02xND6op
LqSCdH0YsiEKByfovvVzdNYQCqMrWCkO68EhTL6O4hPepxm6N12GjXWit9+wJFfr
9kaneiCzFOvGiO7bvcbwX/VRiIGyxFS4LM5SYyEjpOhwB/rfJ9bB915XFH1YwI/T
JRIgdmu2jQik2ZNCk+0WH7+qD6VRJcMUQ/3IL7MCsaBVeeeySJ5McUlYGmGbTt8H
UGf0n6nSCy0EtDe49FcK7ABipB18wVktPqvuVynIDUNSXue6TzNots2v8vWgmZWj
68yep9EHjFjQ2wwykxAebEhlp36wo0/bE+LEHhMCDqrwm3EN/sJ9wRsNxqBkjppM
NJaJqc4Y3J3bYjhNGImmONOu/NhRxn7b78zeKP42AyoVXlBLTpt6eqqAcd5BLXFB
FTpdOSDyOHxQ0kJtDPfV1/iWSaOm63h3uakUXYQ++HyWjpFKoytxhRxpXOXf593M
S8PzYu0Q7HCBAo8sxbM1m/HHto9IoOw5XLNfsVC0Dmhf8TrhEqK9YB6MXXLrCb2B
+PRS5IXa9Bmks96v1IRP3nacY/fdyHJkjg5pm16i/PneiXp7iK9oODfVY8zNCdjS
8SXqMBnYC9pe24iQ1jF4D6+Dp0UVAj1568hu5590GpJGStgpviB+bm/N+IFZcnld
Qcx1gwDIttRHooHY+rUgLXcW2rF+7r+5j0XLLQ64Kxawhv3taVuVKoT2JSEJg0CJ
yUxH3gk+ZM9BMI7SGYC4Q5wNT5RHzP/AKFOk4sF275nZFKZHx88D8gc77KFsBEHq
J/KHD6PiNCcKiDobgCuo19Uu+7ax4YZzVDxTYrev5qAx23wW7pkIWdXsGo1G7jGw
oPV6uWx3iOMP0UsRI8IJD2thCbGoCYdD0fEEDrb2qKJuTn6kyPEcVBpSpCLc7+OL
2BCTdS2pOTxIll5qWBH2LA8G1RrqVzBu30EqvA/l2BSMqAKG33BwiRQfmqYEBiu2
MYKR7DcHCMn5JlSCR1dbaM4T8QUV9hFzeunqUPFujf7LD5Yjxy5+RtUS6I6nHiQu
45kgaVaRIqJ3GiEd1KxYZsJk2zQtujVIKMACv08sTdRYHiVu+aC6KB/iMRJmBwxI
UwKKUdNhTpNLFFbMzvgxrpNsYIXZzqlzo0XjaNLIZvlYxwnDX9AKfCU1I2hY+z0x
EUaVYMvm1XQGW6ALOjvVc0ZY/bBY7aUIwZWPoyUL6oY0MxgIW5jgB5nM0QPObQe9
x1THG0Wx9pCg713NlPO0Q56p1hdIM2fFShXuBYXo+RQIZDWolTNLokBfz4sGBIuU
qwq4+641/MLlQlcB3e79fbEtkrkCEspocHUtWwFUW6ppWU5ziZ4lmUoWQ7EL03dh
Ltzhme/7VLY7K5WyjOLCMXHZ6HGFUeaBeGtwYeoRoYx68aUBrFoCqAMNJ8zduUJh
3SZteL8Hr8F3jXe+Y+50e44GX9Pjvwuvlqy6GyoELZFEutGVCN3qPUvxmwJ3jW6x
xKdcrUNbQ9RZxkC06rd/1bkqG90yGNP7DYSEUGh0Svd6uIXzt8Onqip/gSZxDl0L
VwOOdtMJ/8aQw9YGGeACTlf46YVqn8xQquy2ZymGgcdZNg6lv+cgPrfBbLvfjv/R
Tiz6+j0EZfuKhi11H2BI4OaIdBpmsWSkKw585pC9YjFkPJSgd9n1hBp2VDCugQDR
/fnCVoFk4SmYfnithwGs4NZrAY1D778x9VSIrl4uZofOTn2mTaJbvTN5c5ZU/FGk
upXXY0CdtRG5PUrBJgVRwy0lbGtd6pPG7mHAMG4X1Uy/ASDqLW9GHRCMQN1N8V4T
L3atZgOD4p3B/xyb3qcj5SGO64uXeYeGzhzTnSCw0azmFcPdQNFmKo2jgKtLeTxA
PmpMT3phGsgWo6jlIjLoiN6N31YP4Kn5rANkjGEipUrIZ1KfDvcmjh9gcVhPBePF
rbG65HstibgdxBFt8dMQ4cKEcUGooRzThnyn2U0Poucgl0umWXc1gbjTgMBoElHs
kyVv3qbmz7aa7GO5UJVBfX2tQf4wbN8gEoIF1XHBHxsMhN6UV9P9bS1nwNee/77Q
Hq3mZWZQ1o/yoZsbd/Rrqf28+9q4ZGAU3h2qep8Wku+lUiVjjTYS9nloE7yEkWbm
8nozayLI3W1LHu+Y/cqBex3zwzS/GwJFVZa3Ygak3lpJ000vOygo1zcTpk0Hi8Ax
HePxGB7uWtJNQklGjnEJeGCuxmTiYjk/rejIHu4vtsgCm/oglwpChLalwEn8jcQi
U09+elX1EQLpMi7Xu16MRtmgerX0G+sXDniWFW4thzYrYS3/mprI9EOm74Bhnkf8
5waE4NaMrK0SUOzGyE2YjqxPuw0IEY9YM8Ujn83WcNk1bmcik4j/7dUeR9TPMpwC
q4Fuql/Fik2p5BAp78QSTsUnFBdiIS8uksRtmMUR+lAe7MjGpZu4BbxgqPO5btmG
L20f1VXoQTp/nN+45Dewv2Zfj+GboVfFLl5pteqKTBKXu4OH8BF+EtEN/n0UlRHf
XZal3RCnezGpUW/btUpydrxP/duatLK26PfMlayf5DBpp7Vi0p14J5CDajZ+9w5+
P3Rp2wQDy73wRl10ULK1WhwEdV4vig//1v0Wo82iffYz6PjUv7ekT7lmotwwBv7P
qlwqv7gIwrCU4VMD/xtH3xvrXLLuJb+stoAdZAkoG1kKnjVwIeQml48WAIIYrBfn
W+C+k1a3sv9gWr665P+zpKZFEc5qC06kTjjI+1kYObffkNlTyypiaYu1Bvab6xP5
feP2Jv1MK1K9b/AAgWqeNdsXl4moPyjVFYHkxCMDJpcjcO/9dzjGxm6gpw65XDMn
pAQ3H6iKcB9Oi9tk6iSZGHDtZe1VJmgq7N67ZIZUr0ydm1UVRwlE7WliodnroDaa
4QdUwe0r3h2xmI/qiM6aktDbPaZxuZqBDXu0i7VD4mCLVnBe0T0BYV5ODBcaeLAG
HPwrSirK+hFSFirmAVqlNRHP9MlHqOqZ8N/+fOymEdYjgopzy16KVh/wwnzyi74o
9TDpPrCaq0mVG0SvYT4/RAgaO3MgEPtzjcoGDyUTzv4y1+AD2r7EC52P4h/RL2Pi
ICcd9ybWsRzeWF4pKaXV7T/QsHGFK/GTu6SQblgpSdSYNGrK8np5Ntl1xpZGWlwT
WerEkt4cMOnxoh1cdQoiWMGFEWnH4JzAHKj0hQJvyBYNks8bJD5V+Ss1SGPhryZs
zw0utxO1193LjZGneZd4ub1jvoTEB5eXxCpdy0UYxSKMzcbMoafFDJD6utaAy3Um
7EzPtl9efLlHhCNPS9lVT3sgqyVygbMGMuogN5IcO/j6w/Y3SrKHxgzau5UFo8Vu
JYaoomoryqz8CrmC5VN3MuYBNt/cJ7VzZhnA3Maaa1HTPqGk9MOZQr4ztQgtmkOq
4C+qncrwyihS1sjzx4DQNFcvrMMNhAeO6CXbVs8w7aSjeDCwSYYOIlr+Gix//lvQ
ni0ud/7dKHh8EKsR5vQ7SCy7bPModj+TCFwKyI+W7eCEVMN6TTJAGnmkUFZoj6k6
lqiC136gOvja8cw+zB6KK8HvwzSSNO178xy5ZvBlSVsqV6xEv7agRON4lCmmLJi+
n9cSJGWg6dl0XcA2QLXhhka7xcKSrBCocFYO7WtJWvawpFaEN9/NTVMyUJwUYHwd
tLuiPFWvnLSJM44HafcS9zoOfeLEkGsTdg9cWm824U2DwbEAeECB23+cuxQpkjI0
lXmJCvmNpasqcVen3UuQeS6UXOuaQ/7FblwgywmlauQ5nYu66YZj9jsbiSNqCCMv
APDDYLqjOMN2wE2K9ca3VN/ephLN1x3ny58XVBrM/AbKPAB1aCwS3YcdbaA9QxfG
NTC2hmPR3z1+gil2dNow24B35bXGwyzbTXDW8kAzKAZhbj270Zwr1rgJQd7dHRr4
0cYoU88C0vbFjXbhoG7RjtbClF79ahDR1YehWdk+mgjPlPN9s3XvIhLWRiaPxFV3
hxqw+eoa1ANAAEmOvlQ4RsqTLO3oaVsoY/WkyPdK/dl9DDxrC5ezhyBtMzNImHRv
fAi8n4ngAFItq5XpB856dgclwN+zV5ondOLBAnKvOF0w3iyEYnJzjvoVZG2pc/Sx
hMEvbp0KMpjwaFqJ8Cu20PUmTPIpdKak6GqbOiuW68yxyl1T1RRIOMshwq97NtEn
uV5GgDkvZutcPRHW0KwF/2rx1DYh3Ok0K+wX4z2emov2KuAQwyh8yF9YSZhjDKsm
Bo8QQIqDyL7D2q5nz06yqblgfNwfq375yRJ3/M9WJqXi7/qTz0iZ1Ekn8aTh4Xk+
dHqXLvroZ0u/nqsyBhQLhg7V2zkAlPbVPnh4nSxBWQPxWtDTzDTatWQkF15tvy27
NwN4FFvg8sUu6N7Bi44GSzeDsmIu/Pyp5lhjc4lnyRVIlJmh/67jBEl35p/c3h72
8BxGe0094cCNp7wRR3iSijsYLXQhWrWwlXjn/SK2dGe15PS26/puvqQfY5CLLmy8
ehvi3d6j5gNiF3UJAkwi9okskt2Dkwk8X52C8MkoCCKRDXjTJer9KI40FkLeNbii
gx1YT3wtDWob8KrP4Cuj9CDK0umB5L2OOOv1pXIBZW7D6Oh87PBdQe+lSPqPibK1
nSMxqfIY6Sx1MhU0RJFdpH2pxGYSQRRGySObXtZrT61Zgb9qDmFIVfpiAoyP6ggv
BA7QUmqIYu/uYi0r5QWI21fmfyyR9a9XJZoXjdUBLk2B94ri/z/q7m+YPHpnjEDV
wBnVs8miXEW8dv3RBSUeBSqPz0l3/3GiTUPAuI1CgMMVpFc2aHRWd8AP2zmTcPri
QuM2Wij8snGYmhd2xLmiBXWz7c0UrehwgnwztORBEDOigfsCwKvdQRgYV4tSknDG
LgIDxMU9IPIAwM6Nqoi+aUhhrSWWYCgw+RcEsOELP33wn//76qR5gbMowIH/6I3O
T9QppAoH64c2EQ9IOF8B5Ouk3MelEpRJ3A5rf3tfJ857EgY5Uj0nEAVTJOsyJwFD
M9Ofkl2rlxNAazjEtZPz4GG3FglQ61EIKc92WouR17nXQDvwIMxHj58oGma3zFD3
RypSdwYlil0fmiMf5ghmxywRknvdPGmKr6UracDEoQgaUcSO28TIt8J5Iv2e76Oo
XY9NrRfF+EAwtHKxSXA8L/1ZOVjtA/Zj7fjtVD7IRJJSnWjW58rZZy0RK/Eo0/PZ
AfK69msjNqGLIP0z1Hw4rk60ttGCZ6HZzModgElxvDuv6a8yoIJ0tbd0nHxXz89a
gwyMsiRFe9k/tbM14VAYhd6wPIFhv/u8qahSkX6uY3decZc32fGCJrOUT7FCG6k3
plYAPYzegExQIYH7Lsd0oOXptTnXEOo4zapYD7qNC4lszCi68qb9N9A9awKfnIMh
Z84ZWjZeLh/FgLGJHGsk2Ld350zhMHQDhIJhINfGnwlvaUnL2UUf9EzUnQy7U4F2
pKIU/8sjpBsBc6rbJjxcfcCFPJpUNHm3J+61OpIdnbW/Giggzx/gUpPpYhhwFLU8
ZRP8l9MZVy+3AQDCg4poZD7uVsypEemn0o55MYhUAsrf35103GcSSMEG66YzYZC5
/IonTPLi2bhWk09jgp6b+bwUf+TMFdiWt/wtKStxfUdc1rAVNR1HO31xYac/XUvk
6AukssZEb7fFlsAY7CEHnho3uCKnfPwrGUFPtPclRGKtSx5uZttQ14MZmqnTnBYh
8ifoxHDzgPXc1qXCKvWhraJnJD3jOyeusy7vL5KQ4YMapHQkn23OfyMDuciMsb0X
J61kv5mFO1nq1QLNZC8+WKTldGS8+hb4B1TiY0z4U2RxGo5RHlF9qwDP8lzTFptY
saSkKS/9RPVtSAgY8iZuTHZUnn5mhRfqd3Dd8P6VPgkk9lxpxMdc+fHZLObGfBx9
IOcesJmE8CsZMWmWRciRv9rEIujzD5bUwX3piUb9cTrZ16d5JWKkN/eV9SkR+rne
WXVsLpT3kuSgvgYl0PEhdIuA/6Xot53AcLGvWb6SIzLHANiPTie2kwtaPqVILA82
AxEF6dkLBQ4vtsHOkrjJLr8A7Y3K4PtpkSgLdh2y1SkMpLl+tzXEe/+YiseWvTUH
qAUZ4blasqP6KOV9ubl1E60OV9Yltl9VHPq8QhosYfv7ndbO8yPt60iVPmHdBv+Q
4ZVRMu5E1uWfG9d/CpVzpak2ZF91JY7087XoY9Fg581E4/qnN6MDRofnTDY07GEm
hFvejQMdzj4p6IpHmUYQ8El2UZKFpsx7841tiq0x9vmdQJvRtlwgLDnt/iUZ53wh
6hMntgUwCOGYsPoZfv0PfAarUjjwJJLqgcSInv0ft5jemDY1G+5YoohzrQU/16oX
5hhyPhBqPwt62U1b/NvPHUZCEb+Hse9PG3PW2ec2d8KuddA7NB4EwM6SdLCs14a3
/flkdRGb8qLhB727fxzi7lzkrKCeW5ZPRwJy1QY9Rx7o3NmR99imxI5JkBh0N9Um
oYyxcZbk58LPpLz+t1ajQ9+Qc8Pqv7TLngy215Aau8AII8gaZyNvAC66G9QCzunI
kXqFHMTIr/uXxXjH/IcxRgh/K0RP/8nalG5iIixlyGw9wWEJr6ECf1LqG5GH0yvU
vSEatJfLXh/8HTQk3LWic9pSaXi2y/ZtGIhs1TWQZv/1FCyiehGtQACs7qv7/l03
AZxQXnms7iJwCzOIzE+2rdJGU7BbiF7nzUqe4rtfTVwwv0kl27ZAaBYHz4ZVP+Hp
d5OLNU/Gev5F4ylKLrxAeZNdbMZE+Gnewp4EtgSEssdh8vj6SRKL4BHTfq7ECTea
dH0so3k8GsvQwkVVMLEh2sTALGfpFZ5QNAnjVQsQ2qbbc5GNR7sIcbb5moBu6jjE
dIrT87Sl6836vSgk0U2HLiKux62Uidt8YE85gvi345MvRkaoAH5CH4wNMQpovbSW
OoKIW5Cd20gmJYyvx70iqxdF4riiZcrHWGxSJwzzYp5LI99FABhsam129tfRaTzU
OrdqtP15PNGxsmH5y9vvzCTt+1PIRCUPuDj1oBJzO0SW1JR1VlYfCzjE6agU0kar
T7QS1SK/8pzU5MG06Fx0td7gLJ02IHlZVk7g/NsbF77nsz9zzwppdIx7krO7un08
okI0R/SkSdhUQyFNs8fThML4O52FGSmAuAL8v8UJWmlrPF/FmhIiEN+82qP8FURM
Q4HZtGrV4Jp9JpRZ+3XoBDETyyitbh/SEqwR+fPaFyhFIkO+3KF83N6bCYm56a92
huWMg+RNqfxG0tqQ7qcwGL1Br9Tg6VuiJBO4qsiGjbSz3+ID0HP1QCPjZsyUe34W
1h1g+q+Ykk9Yw1y1RzihvmYJ9XLM9mdLhdsLZblDuxL0pcyNCA7fgLQJ/eZiOfiS
Pzm5MqWzxqL9u82v7f356LPgJeVgrkh3QRdB862sWjtOv9NFHWCm/na55IoT/8Pr
JIKAsa5UFYguaiEcwpZma2MtBNIKQwcQnZgxCLIA1PBWxmr0xmcJjiM0ls43UkfT
YPOchzrdOicEGule6/sHVS4KhlURV/2+AqU50re8ZbxrSc2aClZ9P0XcPxKi0z3G
GPK2hTl5/aul6uEv1cm9hidQpVSAvNq2KoNKVdpL7E4VvN9Xayev6E+SQD+jFcCq
1y4NiIf1YdETramAw3wSBIyvZDOltWHuSUdw8/ovysytYrxFxEE/+28BlRFh5X0G
rcnT4K9e8aAUfAAZJ/tgJ8XcZs7LzxBNmfnlJcdat7a2xV6x+xnOWzf63TAK/ypc
CHAPO2RK7M51q+KBmtkbOg4Qt21Iq1dQu5ytP+xh+7KcZFL19Vu1gK3VBTDd0jgG
7qBgdNpOsPgKcTdXfrDw8uS/dttYTHGkHwNkzQVAdflZwPa5HuGXSjZImcbcd3Hm
Z8QnvzoBmPXPBSuiRewGPMhjcXlCoEpRoFK29romDEDoajixsgyR+1qY066OEov7
e233u2qvOdxc9sYvIBXfNag3wEaGFSWkt2NfT+B/R7EwSbXMevZNN8cnLsbp5SPB
vDK2C+qYvH61ZSUfPCV++G4+SASbL1Nge2A8C9eGac+2O262k5yn4Ydiq61tsCsf
hWG136imF+N3c3KYU1KvZGfFO3MzYpiCGpOkKEf/+d5AZy5tOeJFupe7wltdYtPl
imke4SYtfXSLfP6bGib1WAFXMze1m/5ymHHMQQlEH75YrMdJWK3SwbR5NwWJ2snz
gSrbC8ERhyJHaR8BE5HxIpztw87YFbp0X5gVOFL0SqF4WOZOC3NGPts31wdwu0+Q
PHSCpEbmk9FitjIksn5C8k7yffuwLMlYWIq26Eg8KY1j4gsr8BBCbKS84kQaiS01
6Uhu+gwv8Ph8oZgiOE0KQV7sn9GmIg+pJaCFXTi23BWtM2rCJAWFpHo4MHUzkrn/
T4yU/Thfim+uf7RQkPJqrfjZL8UA2BPE7Xf4brUbMMBlGXkmAJriTu3oqwW4yKir
3VEHS13URldnlQFch9zeElSfJwQuoyFHxGIMhu86leqbMefgJZf3keaHENu242Ei
bpLiBQnSn+TIoHvUTi16PfUYxzkMKF9E13mbCLnMhb5tluXtfTh1KDxp29CLkFzZ
UoR37TSgFBn+I4AfEfdcK4D3y7dsORkY1p82zLyhBhRNcC3bxswqBK8IscE5jleo
Dz8EDi1hOKXL9LDzwZXlBsjVklkK+Jbo22TiAP+gfxdjviEbEio13cR2liAEynvy
HRRJ08MrfSKYIFQpmDBLCfk6NG6AcFLZj7LYr4GNa0Kd2xLNjjNihWSJzVxAOXml
TgJTAQcoILvGiBJqJD1U8AyJ3BgW/a0sSPvnFK7yxjiSeXYDr+Q6gVpQ2lTHUT2y
V5eYz3OGC8kIb+6U1X+9l7ishWMScSolZxamHEL04So0swMLSfBp9oL8rKlXp4lW
NaK6mgtNbAix8idxJFVg05pe5b5DvLI5PZ3cS1Dqw51oBZyeHl4C5mzSPC6rBsn/
4Lz3+U6kfazS7V0Z2TYQl1OGtcXtcVBU18dqNRKm3ML8Bx4ZYI/6ac+qgyDViJbA
RSfkQlcXe4XJfcnSZbCf7ULXK10egoPmzh+b3LGwCRK9wgFccEsF5iVZrm9MhvSO
xcVD3HLlaNPoUEc99mluGEy6u4k3kcB1EswqUniFGW7spAEZTQdRmt9Tvk6CRyEM
F1+7Gi9J0H0r1lqDrmmmu+3fTCYJEivuOapxHQaFGjHHAai4S5NsBqKpKNMHp0In
Y+AlxN/A1kUm8E7VUkdkiCPpD1LHQ8f6U+gUbWsnUJb1GFdh1y+4lCBN82NI1OFh
Lyz3wGIEJWmHIaEM/fA58cNEGCRzrClYx92uANUN9HJwP9LFZgOXEPDhQ4VyPz0q
3a/vQlITEMLFNdpe7DaNDnutsQbl2c6XWl6ZrvLsYYPD5StXd2InMmjtkBjQDojX
y1V+IGpXMg20nTs5lWmnJ3wVvcPUISrvG2aamxFr0mLXvuAE/A1qDCWXhROTPSmF
xBvG+VEP6a3VKtmVRbNX+wqSv/g3skmM1XWl1obZLxJwKb0UxqrPBvuomz4fRzHZ
AptOXHCCXXuO7bIy/2psx39FmzauB6kEUMyjS5tAHER2WitRwKyB3zxTQFQ/w/JZ
WxjEmRpiO2sYXpnJo66DmOB0ZU2FSBkg9VTtk6IhLFp9+kExBpC0Zmgy8mY7O36f
vVa5UE3DvbEthnzBAMTu5iMgBCaz3kFsrTpiMybgI1l4dKYAccCMh6AybD2QuNFl
ruVdBGF/sbUHxOkRuNXHVhn7mdlmZWm55CqkoL6zyAftWbHYsFVtwbMFznO7NIcj
MPK+gVYmkOGdzDlmS+0RNEBkfKezPA+wOdr2l3Jn/liB2JG1weNPxkGsRfSPS3Z5
y5gVZr9cYb8jWo3iA1dizdTZ+LSFCvxbfdIkJYY3yR6spXcNyR5Qjr8eYajvl66M
kBFNwJVCz7qQyV9MQIBrLnLv9CkDggF5GgaXjBhwbS53i5kNLKgVJb2NYi58zwJ6
MnIy4cF8nI1JpbraMKa3bzQdlYyU8fPnIRWv3e9i2aANZih3k+aay8o58bzJ+9cs
nSmGz9iG5tTAspyK0B+nZ0awhI2fg/hSuqKw4zT3xzPdOYTrqG9tTXiFhlAQ0cmY
0v9/lf6ysE4yI17yRXZ216iO+d3fY3HYXh5SmafmEsgDI8/JzmAst/yblMgWRNrU
tE/3jgpcQUULJjxJlF4hAG2bjcpf3/Bdmta546YKD6AngpY4TtzH9T0QUoUGIdmd
3I7WDkfhCsbbCpeE/EMH6arDbEMJ46BwWH2mDmQnS6owxzthhsIETmnCYwqYTBdp
BLTID763yk7mU8dNzvfOd3rVfyZ6VS4WPsz7dPRKtrIys8TOpQHjx1dGVTnQ5mOL
iVEz0XU9bgM3EIF9QjFgtisStFZ2X/cHF9RWjee2pGRvtPD7dZZcuYynsLCVn8ji
hrm+94wLwK795uW2SuNnOBvjuzP6XsEaZevlswym2GEPBGNjOu3l2WrZgL4Ou0kG
MG/QYXw8y1H8TtQtgBbIbgLAca8Bx9vuY1Oc/msH1ROCN+AuBzMq94PEbzzEzkqu
T0IjyCIfsn6BbeZ4Szr6W9hM2tM87gIuHE9IpsGnqXXM/RZNGk7Yr6jTpshP44cv
NJ0nkfCPbhN6O4L57KbyDqt39amyvSQ5Te6U6h7k3vcvvhCrFxPwo7sdsp+6Xn/2
AueDtpWuhhwNM4jOleGz0189Z6c649f48XlDCcNoc/QxxHMZ36NCskm1I7+dP1ar
s8Qbk7Q8MI4votfz4QtKI+VjZxlherujHb8cngHPQ9Scp1je79iCOovZp/NgMJmV
nj1/r0X8vs85vjXJRhqoOpvcYY5Q9R2a0oV9t3IzMMfeLlsivl0+QKRBbBkUmnb5
ybuINMrqBgKYlmabPuQDOTyWg9m1BcpHmLWdv4LEEbFQ9y34ivA+m84PUylit6KU
+bBBNIa09n0RtsKXz99YVrIJ/YY7wN/fXDHnmv9eVSYy7A9TeYW1nEI9r2qEQHjv
S18Xv/Uyt/6FS2Ylirt43+tt+sFP78SAMlvTuWE4bPoLaYmx7xqSwWf7OWY9HBa5
cYEieielgoV60JQoAfswa8zIsvPxNkfahlFA1OmAAJMo1CrvUw7NGCWQcG7HX/SJ
B7MAacmIMiKXinIe7ptOmi6cFeNRVdcHY9xUzTyWbSrV+9OWHyO+sW+xvwePcuH1
8v62oQHg3Yeu5RenkKh2kFxTHQ8eZqBQwT8F45nD0zppLMT5/BqToF74+MU4Vtfh
KbRRBxkAkAvVhnQOeZwAyXS1c6gLIoAcUaz3kipgF+OdAUPwUGrJxZI9daRCNZtB
QuYeB3iNBJP6ckf3JISJDqV5tlpV7NuLfnqxfJ6akY1PdT/BMloum9FWV0yoJEOA
G+5N01aS8+zAxtG2gF8vfwnBCFYwtiMHA2q2onTzJI6LmIrkCdkKadXErjshUyZM
cdN8RF0x1hF7KHY47rzZBXOgP7PYMRFK8Es+mhUNRuk/PFhRLes3sFLPSH+lErRM
uN/G0VocBzSsLNuGutWFRwspe/Zimm6SMd3cZD5xW5uV9uxMwViVUV8pq/peKs8L
dZmkwPjmFNiZGkHuYJdmH0VFHWVP9c7H3eiHLju6Td6mU+Oe9gtm8yeAPrTh5Vvv
LNiPw0d5m6Hh0Wlft507GAMkBDjsv5qUz0cQE20UPZQYr4fu7XDEqhrn8xwtp4BO
WsILh8a7gokk3rycWPnzwa5pLBsXqKdFDGN71TLky+2mx8hmFvBz8enSPtP7+Gsw
cCgFQYUGu5P5DBgTD8yE4pdG3t7EV9Ora1Q314WvB6EeUnyexveHAM3LEHYfB5VA
AE58x4UElAf4EzJWmM3snxgmQvTLAXc7E9B8P49ZioY/dtlioiwDhga/4CP8JTIB
DzEFmT5jNygc2iR3O2j2PN+pU+uYgjqu+isKiDXo9ztGHATUfvT9VqM/hktAIFEJ
4uGZHp2AFPHN8WWKLvuXhk9qVIOpisYiexq6u/1UUl4+lzJl3uXgWJavnaPTphPU
RoJYWGeoHDZHTuSHj7M1H5sekf6wL6jbDhJfile7KzkifhNtGdAM99kx+VMMUwsY
Oo45VmA9DS5CFqIAVkEcDcFh9Op3iDF9wF1LoDyVURyVIxjGsb4UUflCXmqlqaD6
lgXEs3VXHIsyqn5v3JP/oy/SB0sKYxdrv7vpmXL9AT18Cm6ZbjdYsqcEoI8Vc9Tc
lfbp/Us3yfuEJ25B5VpZs+6Cryv7HdmsafG59+DPtiAj99By85SB50ODtn+jrRCc
j0P/qu7hTqs9pY5cp0q5mnl8LRbG3dlqg8jJKuImKvi5kN4oQl2cozP1LsoDj20j
zOG/fJcS8FghPZ4gNon5yQ140e04/N3Lf3KdD5rv/1RG+8DawmyUhUNI2npcZEx+
kQPT2i5waXBmC8kZA5jXnfoH+h9piJtkf2HqqzuYf1yQAP/MWbd4Z1UKDjBUKZmn
Sqn3Z+NdxVlmrCNuAwSCVkjEaUqel9GvM1YnC2tUdK0DLQSvsh8KiqFLNeboaWOO
8iEYO4uFKLsbjaYRTumEaWJ6gY5t3xhaazLqYqiCHuAmHNV/OKwOA6tfIPZodaBQ
jt59YnYVPvUYSxZLt9mG1AoVcgIT1oar/ARaa7DNfP6wDJOj3bDEKF5XDokRnxrd
WGsKTlJ0zfA6hLkun3oLnc2suAO4Bj6fFkdZwBOYSst0yf/neGVqGdMlqWZPiVnk
artQ9DKt60CAWDHJ4jRm+bTBCVCFB/kU60pW5s7Zq0N7Zf95+eZj9WqhV1TZv8Zr
xufB3OZTbuqNcUsl3J/wMhoQ6adopSrJwkz0qkVUGc8tVaf6GuRscl8SGzEcIbGZ
sQbvbzaaf6skGN5MnGnL8+ENTnvWna+pjc8ba4mYdTLl7u0QX8rfViE+5tGjAD/J
jo4wb4iuc/O4axziub4zD4115yZIZzzLSmy/GFF81TBv5wilqgFaucurcQPGT2Gx
FKJ5ObF7L1vS8NzPemRmI2abnB58Q5FBN1vLIhx3iqMgDuIqfXoZum6kaNrG2xbc
tFGQkdVEswcSwCRWcpGOobUIoobzg6pjiAptdhvKkKhYoibpoAmPw+tClQdsAuhF
J9122dfFmxZxmC0IFuMdv2Mf7D6vzRYtq2lPZUjpJDnOUlWZoTuxq6NoKeNePNNP
4t2dcHNv+vhPjtIBqucZG/bKeQPUsrKWBpCCjVzqsQgrFhxAbQTowWZ3tUfEAwnP
ncpDLpS+RDNG5iHU7HnFyWLVCCc+F5qPz03CcOTeGv183oRY2DAsv0kd8pOn9Dol
Mb2fHQyeV/JNkBaAzXmGCFUqrjiq76zo9ymfozZFZx2ud7/v28AKxj9vadkpUhWJ
PL2UlGQf734X/7lnGIAEMaCRsyjtNw51Y2XWTr2U2tl1cwCx5p/QdRARfb6kQdje
dU/316qw5LMmLFf4MSMztP7h8jt4dSgiEgk/CpgkQEoCXJ2ZnF7gugcCdytsg3T6
BYlxaks5t+HMQyRuLa9rSgl1Lk/lSSjj3oqDiPFwnsp8SVumSjk0dItTiJQuK3xN
bSjb+AnPfwSNu9DQXORNvBupIl+PvlE2+FHTaYSLoAUbIiv+mWtwnoFV/f+aUXqT
me3ng5um4y80aRYnDvnma7hBqoqH0AVvfM3JBPmqr4+diT/lrZAHQ8hccF/jv+MC
LzfS838X6tLgRSpnADy5mYWJHe2xwfp4Ee2R/RK+A5VprQeKFs86ud6fhjicwVHJ
4pt4Syb6bqwTpMe/27YAGIvsZDFv3hX5P6JI5+x52zbNqn+hFs9JGJobT+AMGXgv
/icwyvtB4vEWrIqlTxoVVpavf/mSqGz3wRry5fGNCPfmbbRrRLgr9dGp3nThR6Ec
L0C7TPF7hMNsYe4e14tVnDZh2H09SfxxATPkwVIOqfx9uGX+Hz9GTOOzdKzR1DP8
OCDx1jT63eZpyJAJADcmgsxx6y3DraAWV73oVSDLjEGw1fXFej8ITqBT//ThWcA1
egM4wGziHpOSzaMgkzEk0ORG62o0ArcDbEwfqtg/g+fbS3NLpdqIQO0Mrcxgpld+
e9/9rtFO+B3bIIEzxnCFBXBc0+oUCNQi4pwvxYvjLTtbFzuIbFbAOA2wJjexyBDC
ahYnZ2FQVrVhADosCshsbHr8XHWiDAYUAs9BP2mpsZmupi7T1LRakRQDIbX3uiny
95P3FPKmDdZTsgbiPdKnFVT0cTo89jbu4uyXeAoJJ3P0rV0of9/OwAb4OmX3mzXP
KXHC41U8kRykvKbw9N/fkCN3QUzQuNWsQ7nIoKzJ2xVqj7l9gjSubTVEXzSBIJTo
YC9obhERvZLgA+aCSWGiltjlNSVwp2LO7/mCb0i46ML2qhqy1ebPZqefbeTeFzZs
TSS9ANmJ9kcLRwmoChu3V+JSyf6622RUblkJ8bCFRKPMQ1IHzxJWmZHLt7Hw8Cuf
lOIfGEktycjDGwvF3OtDXDGMFdz92uujKgRW/n2/ihtImtdgWZy4NjuFmNuZmZ46
FSJACaUMVnYis4/acYCm4ElzNMozvnistDmANpMow1b5mg0DroPlhEY/qh6ayYeo
swq903NeaIbgmSFEtFfpwspoQV7TXsjT32GrCZu6cwL9C0VJetQGyxNAh75A5rsA
p4D2K/z3z9yO+MR0EdumcZkhei4VQ8pX6poEKdAGl4CjtcnsG1/N8ml/ns44F9ea
32bAhVahJrGQgFgGJUEt0v+1BpMITnoF+0ZCKssMczb4pkZgcIgUPSZAyEGbX4I0
+2Hh8sFa+PiyPDsM2K774cR3um2E9sRCMrKKeXzZsomGpzSawWbMM/oTju7AMwfn
bcYXG/Xu0o+39PnTOid0c8K6C1qiGq21RUyQAo4AFIoehRwY3HFhlDPswwHlqkCJ
aWN5qdazbqMSSi1W4r1aL0thjCS9mJZdB0CpT2dn3m+KDrv5Cfr46cDZVCYAL80n
9WzZ6CCaOMDZSJ//B3mO/pImm7Y2VdITQX04sRsKJCikDPOYjR87IHYvf9Kh2XDk
RvGIQpnNEbKqWxv3/PIkT3Pt9NUMEaLMNv7zN6Q1WOG3102x3yTpWdZcga3rV5Ne
aQ9dohZMW5bB9QhUYwhIaGubsjJh2jtoW9LQJUZjyhDzNZhZNr3rC+w/9751qxL/
BWeP9x4yrKKqjamF+PmyPCjPCwWHp135N7AxxZcmhC1Nb7cPRrj3gZSnPMPxJVpV
RToF4jB+hQle9EQDq60o/aGrwngMS+OPLw7QWtGo6XCVT6g94TtjwCTzsm6hnuPd
YLmPHtIWP0WkwGQgTZdB4HGkv5vKozKZDYyunZMWHfwybaeFKOHRl3ogjU+Hvnei
M/1TehByTjjQckVVUR9vwWeyHtyltkZayyEn0J+fT/jlzv4OtR4jYmK+AtR/JWlb
yDUeQ9CtJGWoejcBXH+eT5Ly/sdUl0Zu87WgLcX4/NJN2EAcBDxZuf0ydTkuFjLD
/EPWgxx5DR7ufdvpHthRERS0Ky/zklMh60xBs7s60BRMLzPJkvWfYbOwCib2DMv3
VpOzjqh9oDeLI8WV0GwGZ3DJxH/+eaWjigzdbqVzfzFktSoAvmIwyyKX37TYhWUd
iq2m4AzpOU1zhXUi+gzx4ixClfb+jTBvAtJ3rvOmaUbu+a99pvuEP2Z2gtbdZh2Y
cp4zgd2gKlCZ3yUgzng06Di61zqOk+hxhBPz8IP7eCPgLfq5f1Xi1S2x3cpPDmCU
GJPrxnTVStG0CuiRn9Z8cQ/e+h3pDq9+vtJsQlq7YhM+TMtPepUSChQLPBt4sOrD
LkwDrvIAfiwUW0YKws5Oavf71nAYivJn8iG3td7YkAu58ekS7rWC5+i7OA58z1Vu
XzsMdOYDvQRnu/0sEVXW39Lln9UK+zsKx0XF70yQoXmiz+XHhJATyGS61bwQVDx/
E1lXkrX9Eqtq8wSx/0eg6PaVLI843uZ6IzD4oY9yepWnF+jmMRfyOa1Q7e9FBj/N
6ahA4hdS3jW+Eu+E+6JIGMXMw4gHZ2lBs7LWq6TeHoRQ2ElJIJaaN+Z+Gs2cqmOT
n7W820zmdblqtOEAs0NDC1lna7JIkmshdDAEE9PmA3IyAafTeqiaAYHI1LCBSqH+
tetg3+yL+dIxPyMLg25Iu33vZlAqjDftudAjLTIi2dm6gusZ4InyouNIUS0UVuw8
mHG7F7GdFdgR+krxq+K8vFC92KLsTYB6yKbKs99Q3ovvFs/+NXlPQkkcWVuMRjLT
WeV/Zu6fTa0MCMrCPzU641geojr6nKIEM5lWXoF8g8N3zfNjju5TJahmLEatBmgt
5Cl0w3lgm9VXYKyCK8SoSnOEZ4SC9jxb0g02JO5CY7JIjWdPHuQk0/G62DWAJBX0
Sj79pnGr6K4MvG5quiPbcImulUEXxBYxon5/8qsJF82rtkByQmhJm4pmnGcOLxi9
Wybe89o5yWbCGJVPLvwzWdcc398iIBKEBOkVD+nTZsHuY0/Db0WF0c+4KcrzGbNN
CFZRFabduyq4proPksmeD31+mhqMLAi7BjWtVLpXj3lcLpJKu6ZikF1qPh7Qk1GC
JdVTDr807N7IoyLjZSZiXv+g8W9G7p5Ma6qkDZQ9De01HPYMkoQkMrxtDHylehpx
ZmlwS+bWwegNcpUWcsX/LENovqCJAjPL3Z3edjNgLN1pbzXYARGEjzswgASB9XpZ
WQIzDMBqlCjRjg0/JaGJ9ipxow/S/4hfZj2VipZPZgDe8PzPsGZUWz0INV7j9l6x
6irFmu78iVhSD0oDK7ouyAwqmwSiNaqEwetc1VbAOyVNTiWMilDyal4TTB7775n9
viXa5JEVPBPqiZkTsHx0IfLQtlnhv5KdQWWgsACDSjxaYdFeo9d4FwxNf5aQJdFV
rSeTwbF2fTIxyg481nscuF7tgI3iAFR6wwvSmfE0EeeGIeT+b/cEM01PbULjvkRd
ZEWCPbhz9z2D3KZtjF1KW+h5qfTKDlppQiamYVEYnG/GpIC3PLs3e7lZZ2RPo649
Efti96NRX7XwC3JULaTUIDWsflusn1lNiQB1yIlxXInBQwowv8GqU4sJAQ9Aj3Uz
9ts79i5o8TVj0VVyq994yHD2qmDNZIIZep9LyVdWaH20ilkn4/Szdn2PPtGuc37m
bcZdRHNn+8mZ4hCP7Pt/OIGfDQ5NXNba/1gBV/t3XDtWOvobpt4nVwtunaWlO1PK
55NVM96eQpoXnC9B5xhzfSIqjBent+aoxtyjJteVnATfBeu6mSjWuh2dtGyjvNDZ
pi/Orm4bH6Haoq/1hzlUYFGj/ZqsHbAJ+Ktyrxnt6ALfPj8qDOIRJHO97BYQRFMq
P4nEWmU++RGj7NxzBb2uvjvit01ECOAkZ89/e7Pewy5Vad+tvYWsbWJtDMiKhWHV
Tjav56GGEgwKzElOBq/8VwfHGCjAsaybKm1wUtCmvVgsiRmLDMvqjOXod8U1h0k/
0gr7R8Hrl0sxDxjHldKrkIKlX69yLbDy1C1mPWQhGXHxCecNBXu3sW7ZsvnpiS6H
`pragma protect end_protected
