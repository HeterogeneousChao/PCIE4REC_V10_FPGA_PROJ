// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:22 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XYMYUuilaxWs5qoHU+eQKPFRegkGDa19B1GW98RGZQyL9OBQkutObKAono/hsbM/
nMAhmdutATI4uIIB/yueUkSU4egDa1rL0HY+WmDv/d+yTPXLcIKqEavHpdgxf7Mm
Qm/CI7ddsEdGPkxBFd4uifypKiz++gHlYcjW4XMiAKg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5216)
avofCrnbQ0YngHEqd9FivbOBIE1KfQIU+lXrVwXRkSjEtFerUt6QCwJTmApm7M0L
xZusNguRh8d0rC4uLEkmYZHLr65G0UTSvflyFjJOptpXI9sgn4AS5RyLYrFUvzIV
jyTDXsd49Y4xgzYhFaYasZYv1IfpSyOajBb3laHIbMWSOG7HDyj4yCPUSQFD5lX4
2NOcw40Uzz6jmR2MiEqVM8HPWDhoYhkohzt7fQZxamExC5imgSuMrHWTsXduDgHq
ORXpzS0JRTDJyGd6YZYkMvyfrn2BsLbR4QbTnvda4r8xFHUUEqUWtGooOk+KBKHh
3DwWUyMIW5upB8NuHuPLtFlNA26A87n3svSjZSbQAgUXhlPpJdzbdV1xn8AKywKX
V7KeP8zwc7HgitoqT3xCDDZvF5QGxi3hDWD/s5BDg9yKPocLtRmATuZ7uwApG1rA
pcteOybLlgKeF1l93jyuN73PHes/2PH06J6U1tJ21PJqQEC+6TFhmVSjES34+T7b
yOT1jsFBI5XtZdgXqAlZg8cS/nVd0WJmWX9tKSUFxeloUJbzgtF1JNt4KiBFv8sN
NQfo6knGYpWIj2yJcVAqIED3rL0fgwi5mZvhHssB//ameA50f1CH8DmLgtW0vjwt
bW9JIkBPN4ZPnGGITMH3XdpJeeQNwGeLVjgvOPwVq5DrBPJk4oTzrMFfS2ZCgwLa
+vdSJuydndBFF7Dy3AHTZJbaltYwT+oG7AW5LDT9u8wt/egPFCxta0bFHPVHcOKu
GUu261BJU1Z6bmLXuML2VZxR3BpL7ANx/gSbV+KY3na/BUOSSvVcXs5XgU6pS9cB
Oi1CJpMkvrvj8Xx/ZI+e5Ot+0O+rAk5IMRbpnhvAgQesj6rViWyAqiumNkrVLMCy
SdifAT65Q4ItPFzaU6itMBRi1LyshQzu/OCTyHqLEwbydZiF2DdYPpHWkzJJdZ+J
P6M8JhyJxnpS2H2vNUQzfBqoJUFWgdIE2jRZZlsmEb9OO7B5kikhREbMIingSERi
3v0xKzu46fVdUbIcbOtf82tOzpRpjb+QiEZ2JOoXjIdmW0ZDDjx7kOOAfjouDoaM
UGrxuXzBJABuyt+/ZU/613WgoDKt8ekCGR4e55E+8EnMwTe7bHPkbko2HYJaSYIg
Egv6v0Xb5wV047k69zenoUc+5EJ/VO6ZrT/RIWA2PvTMzSasa0kDec6qX3fd5pzn
7NyXS3uQX9w4RHPVolpyvXwJAXKm696JkrPiHPw920Wr06tN/yBiDixsQTWTNEjs
JbhYYxEIVZPjV9/AAihSsDyxslAYmZVBKpo2mnjslDew8scw4RQ+S+JkW/o1+c3h
tdrv6NkBE8QivOiMN8eseO8vSiu0Y+VsWDLopoVI0rCF8BDlP357ryrim7wAMtvN
uEdfW3nkTaAxoPmipgSrhTJtep0I5g0nBnNqecEZ5DN/VhXix4BJNuh9XhrrrHSm
FslxjIiMqzJYbpv850t/0LqaUL1UabdUEm8QAUMrzV2vZHsE7EmUnidPPsqCgHok
X4WCsyLnm/TQpV2ydGo/HJMJg50X/W5qh2sOz/7rl7Wn0A89e2uMyzEFP0y7LFrp
FZXw/dms+r4JWkNrnZDuEZaVYZnMoebfy2QkFlDrDk9+jb9RFvYYwbgdaZqUP3H9
WDZBW3bGpOS0/nc4UOrLqx9h5RYknk0mJO3o7Fgf3bcj1ya0SNH2ji/Mbc+qxfXh
okHxWg3hEhNHizG843NuWwhFW3KiJ2a4t2eo4NXn7ZHKC544EQ3ObNgQxLoouxLj
NL5nMFPYvfDLLCEtyKIiA2TSo41BWT6Vp3UQNtGvzMTBHDaOpV0d53ALBrHGfrQj
2U3AvfIRYMjVlHyEWQ1jtkZPK4LfY4YusXKl5FA4IOiysq3sQ4Oz92n28xXhS2qS
Cy30VO7UOKTHEtCdC3Lat9zVUUBoGSkLd+x372CymCBZN1SGQzc3SN1g7XRvxEA5
x8uqTOwZnK0yZLzKvGWGRmG8nvuoywVN1fNWsN3xFS4aVCQbdPz7wHoKRlkPQ5lQ
lrZLyReVuEL3w5sU36SYhYN7uygomvF8O4faIq9emq9j9gXfe7M2gAbpdAJz0oB8
o2cT4L2V0xwNRWhroovT1IWoImKXHnj9DHXkfOBpwWoQqRYqLJViZIDk99GmjcQj
JsxFNzE+Y2NQQcVI48lJUrBuTw28oWw6DJM1mpb1ZADNdklZaCQAh6j3fQSYkZtp
Z7SHFaH2arZCSH+ZZoFMa+S4harH/IRJidJ3Zq1hm4tCnYoSfDDuvO6ALQ4YucHZ
RV4MXFE/DemvLlCgLsqTZiQZKcMDU1tkJRg9R1Y7a/aWtw/UovjiMoT3nbIsxhFU
Z7uM+lb1CHIj0gBSep+cdej/QLa82+7mMo5Owa3tUimdBGZxg+GeKh/cC1DHwP79
g6ErA6S8CyfCv2/n3Z+vAmL2KMsvln743EOu4ziy8d8Jo/x/op3RCBGeiEAzNKHJ
2IvX1OgE4jk2i1QUVLxZOboij84ZDMGigtkSTIhT9UHX9z96y6vDZsAFBO3yqZuF
uYeRrFn62RItEeS4+5HaOBUNyYLu214t+Pz1FAlqO325rGoWR8FIC3XqAYb+Rhtq
wtNrV7XkRa8LyeZmmB3uF2ZiOvZbL+/3UjVco40NUT7VcJhbVnf7A+QuH0l7Lfi6
BaYXgDYu/EZ+f7ydu6NNrp2WOk3231+Zd14wDLFpKCvbjXB5l1k2lxNPa0EPBKYI
J45OhPt6kDeQI4TLPRFoRbOcDdL1EC7jOrId+cIROK6pZpRjdsPxX75pR3fwsIrX
rMRAEztNA+JAKJRyhoLGAAUEqajquhab9a+kKhTvOYK0rpOzAgJ8UMpAWRJIpeBG
JV5ZqiDBLhF5DlfBdP5jdGHqoXrFOKYjGX9w2QGTc30rP1FUEE/BTyCOrCM+KyXp
MiLRcVtzg2kVino8kXEPfEtdZ1WbPEakQFFPlqgU31R0UREQUo7MjWgibclGn7Yq
9iFYAVrUOn5GTp92Kb3dmhGIOG5p+S4uEVahbyt25zpbDJHBSYvwSugF/sHP1wj8
ZSBi7I13k3I/E71J39xVqBCjdxun1mCQbAXlGjsgI2Gmz7E2tprnpR18YT20UMWt
Abd3DIFZnouvvcHr7XIeQPun4DHxMWtriqwLlHG9YzDiwhjL7tZthpIGG/YtVpgI
/FZgqlk+4gX7v3uF1m0FAVp1teQvTYEFcyqQBL/Yc4Vr52CdaeDO+m97lVvC6PkZ
yhzXxs+Fh4w8P2G7GBPk0VOoSa1I+HdkInW8sT309QEnO7F3FFHNFx2QeageMrwE
ZRwQhVt+fTrdqFWx3Zh4T33x3qOa3Wjh4jCf5+g0xts0jnDs05T9cukIWQntB1nm
Rftx6o9538DCGRx9KhrHRgY669+45yF3hQhZxruYN5n/Lsr+VZBJNQqf6WswN1OZ
5hOA2MWgXMms0VOaS8nuNRbxWMtbEdbxWTqCl7QpKJV8sToQCte1sdOT77FMDEB/
vtjVPM0F//i7pdwffU5xI4kk+kZyZ1YPhsdNzkYeW2EtCZDVVvCzvZWipuIsD78q
Tb6tPvrWaWphYmAV9GW6IRAbJ+MdXOdK4R/Jy7jru35P/PBsudOVeEkHFKpJRgNx
RbmktJUY9Atn7aiRu4d5kuWxxHw1wzwlxBws1MkTThDbDINhcytJhX1AwT4G6/n0
eG6gE7uKmjQ1YYkg5+d5a35YrJKmmua/fHJZ6yqrNhKhtOqEN4FiLt3pWghrT/Rb
lTb2Gey9XmQc8oaPyn2L5mE1pGDnFvsYuOK2rPdeFpcNVr7JgmVVoilOlhOy/hKo
KzaJe87F80o5Mn1YRqXwgxHg5VV80OzrH/KrmdLuHT+wwKPIUs8EipNzYUIAdAJ6
ptQ7428gp8wJF84BKsNka4ssaIIryOgUVsLiyNPr6QH/tBsbbZZBekXw+JhgW5NZ
CMsh84L1wavP3b34ifVes3rQhuuGUctV4WNFlte9A4cJLW1MdSCQeQ4ZnMYkxomh
yEOlN+AyAGW+Lv063AFUVr3QvX0e0Xbc2rQ8vw/8FxYKIk7F6vTw/ulaxCVj1UQr
LYz3UC0hoUjXwW3RIsod6/wzfT2KbITwvB+1fNrkW4tNVau08tZeC+yVwMEvxmm8
2MYbcN/jZ8a75o0TrKUEXnUnrsUoev0APNoZdHwLMZ0uOzxhEzFaSwH/3FjA8Tuw
770RZxB1fAMMJjCrJ9HhEoPGxsPDJYilcq2jGuXxvPMehdRs51Z1v8Ma8S4EOfnR
JhHlrPLNmfZGazq4yFLU/wC60IO/voigMHkYLA3TdlORK7vplVcHrzp7DPoMS5kh
nGYnbwiMrCK0K8ioqxmliJhEDCj04Waep7toT8yL4Til2+X/eBp3Bh9cQ1sR7Iqt
Z6MuSE3PHI+c8we/KywrHQYuwu0Oh2wgaEFsOqCuJAh0cCiBtdsXUhCBU2V/EixR
XxdN8hK7SWt2S1kxUd9BO1fiKFbqZKA4l723SxAYdFTXalT8mnpuOn5s1E4hYp3T
C5f7kFSt3zN6r8NvXvLBjlckCQlU7od1HgAZoMfUAHk2pPXR7EjcusdhNOcM0Jzf
zD0s8mPHqUmIj2LGX+sPluk7XbBKW3psZAhEuk26BoCp+v8KxEIs1WVESaEJoEtd
Vp6lt2cqxNaCYknronyDWtz96KisNW9vUkNRgZHgm5iDsCp5Q1xbgxVbZQVpud8L
QT2aeBqT2FyBqM2vJOlrnKs9zecevHno/MpehFK2BWr2lBHWcdA+uATmlKm/cI4H
cmKR0xRosrg+GPJ59U+45H2tphrBw0Pd0is4MyZxtTxVDAl3lT8BibjJ8h+cd9Dq
T/7EbDb4hCvQp1dmBAtq856VjKMe9xx0stl4U8YLG6LuRzF9ftmwz/Uj59XX7nJ/
2dNLxJftss7BaC0V5IacT89xPAokHDjhD+P1OxtNUczj4y1Xrts+FWYcW7mU+8TV
SEzdnQDmwMnpG9/3Cd/VQLvw+YWkXchYrDLrmC6rt13qNWJqvGAf5dw9imh2b28B
J1/H7zVBAUTQnWczN6mBxG7oNRjYfU3PtUjNBBdrpD3iLYgqzNTknGiXQ+nV06Et
pOVPUauSqd9CvQC9zj88CFWBD5OIk+ZtIIOJvnW4CZYd05CYsionmQfBWOSYv5YJ
SpfTjiyqrWHmcVuW7XgKPr5xXnaHRelHaVVP2IHsLBK0fE0Wb4J9/Ncb8Iv2lDvY
bcKqy5mk92FBeVakgihCuUnNApvwYhj5cqjpQcs5xapq5o61JBEt1CHG+suVCrEW
jyO3l9PmfjHa0N6c/99HWWma2W/nfjJkwQBQKiAcv7BEXei3RYufYiHLcco8s+9V
0Vs53pE/bacE3WQmWN9Pq2jBDx5hfpOlTPX3Yr7qmmAvnRjKs6ukoyMfQ0WyEj53
7ilFsy5bIdIwxe6mQh8hgz93vU9J86aRF8FHRotWRVrw96yZ3BAgU2K+eOWtLvGj
T4afr14cgaENoOJYSHd00Zwxs7E7BQB3C861ZazQYqZdAdDDUtZOCOJYudkw0IsC
k1ZdOECoNANlGdUHPdFalqw2xyEI7WHgyM7VUi2SVBafApNKg97skLTqo/RyC3N7
alV1E+Qtd6uiLK6wZZPuunnFkTPcf8SVtU7xlDhrxm9OL4V3PvgZC0Dc7OXryoq6
NCaEF412UWB2yKCDmMzHKzgecPkxyR1+rPoJCmNGC0JXuehvDTTnUcjWFdUNxzWs
6K5itYToP7lfTxH5v8Blkq21C52GR8qbD3acg1OXAgF/TMCdb/C/6aBLPK07RvnD
RyAreW0aelfmDh0rJnQfyTYYy+f6C49InlJwwIJp0H2zVkpujt8zfilxR63vw8P4
k0zgYGo8Go/zABPIQzrDQ363h4VFoF3LlYKAry70YAMARlKkAOVrLKYD4mk/ze9u
FUNxFyTKlsCVrr1iHilJ8peIndrnvZv3DB5kUWCrVmo0Osf6aLlmTLQiKAz2RGz2
7FoFxAHnX8GCIvAOKr1rsN6qf2eVhOOPT04rbcAinz4THJZl47oycgWDHEtBz+fy
pehOqG8oqrae2alJgFZGIwWCzT03SQS87TU0JbGM2W3LNRxrbbh1pjX7EFR1Vy+a
THVUFXc/05oxPvf6Xsy/dM/vEafHvFRZPOtyAKyzGqZZPt+uVkbbDxQJvHUqckmw
0BDMsZQnutx3BwZiVOifPNtCExLV94tioEvvPTqOTnt/VdeVcHG3nyRKBrrjoXr2
OofX6vE3C766Lxqgcfr4Cr0338332EchDJVK1k5DJD9J9sJkV8gq4vp7SdrZmI9A
e31NZbC7aVRT/Rd2RMh32rhXwmofmUXnsGPj4ZvPweXYr1CIot3TE9TUuLHWlLO8
7cAFVeS1xGPAjEGKO9BQnZj7jiNhAGbfFviznG30rqigx5Kw2kf4vtXsSL+aaH43
zmM6I2X3I5snsjJM0MfcL4KEhlU4aesxIcB5/6XwKaj9tU58By6afWBA0vjmpy4P
7wvJfCN3c1n0DnjNtO2emkhC6BcFNfnyUGw8kqMoEh3ClfBZjBfeZ0zk+y4Jv87p
qgRwuTguZjlskU1iopwkuBBguraY9SiEJT5L1xNK7CDPdBj36pDUVT2Nm6g2bu3u
kmNNnu1j2157y7mKLcoKn5OQK6A2SQ6b8cTLR9xgbCjjFnfaGgi0hAI+W7+mAzo9
zEPKt2WrAqM2HGSi4UNLpF7BJZ3GouCWzTLFAst0O4lxWQ+irR4sTVBbRdzkVE4N
+waC+dG57vq+B/W8OljnyxZ6tJOT3ISVaQmAy+SnjHLZXt4Vs2HOIf0JvDZy4Kfs
3FolthKVcRIou8K1ry+Y4G4xhrAj5nVCK/5QOuW345QvLtq3fa8s8jXngoX5928i
JP0aZ2ryG4vsLU0+/EuxP9pVr3l4BjbV8zGK6l+fsvM=
`pragma protect end_protected
