// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 15.0.0 Build 145 04/22/2015 SJ Full Version"

// DATE "12/06/2017 05:21:30"

// 
// Device: Altera 5CGXFC7C7F23C8 Package FBGA484
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module RECONFIGURE_IP (
	reconfig_busy,
	mgmt_clk_clk,
	mgmt_rst_reset,
	reconfig_mgmt_address,
	reconfig_mgmt_read,
	reconfig_mgmt_readdata,
	reconfig_mgmt_waitrequest,
	reconfig_mgmt_write,
	reconfig_mgmt_writedata,
	reconfig_mif_address,
	reconfig_mif_read,
	reconfig_mif_readdata,
	reconfig_mif_waitrequest,
	reconfig_to_xcvr,
	reconfig_from_xcvr)/* synthesis synthesis_greybox=0 */;
output 	reconfig_busy;
input 	mgmt_clk_clk;
input 	mgmt_rst_reset;
input 	[6:0] reconfig_mgmt_address;
input 	reconfig_mgmt_read;
output 	[31:0] reconfig_mgmt_readdata;
output 	reconfig_mgmt_waitrequest;
input 	reconfig_mgmt_write;
input 	[31:0] reconfig_mgmt_writedata;
output 	[31:0] reconfig_mif_address;
output 	reconfig_mif_read;
input 	[15:0] reconfig_mif_readdata;
input 	reconfig_mif_waitrequest;
output 	[139:0] reconfig_to_xcvr;
input 	[91:0] reconfig_from_xcvr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[0]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[1]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[2]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[3]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[4]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[5]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[6]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[7]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[8]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[9]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[10]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[11]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[12]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[13]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[14]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[15]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[16]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[17]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[18]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[19]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[20]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[21]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[22]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[23]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[24]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[25]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[26]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[27]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[28]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[29]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[30]~q ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[31]~q ;
wire \rtl~162_combout ;
wire \reconfigure_ip_inst|cal_seq|reconfig_busy~q ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][0]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][1]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][2]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][3]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][4]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][5]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][6]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][7]~combout ;
wire \reconfigure_ip_inst|reconfig_mgmt_readdata[8]~3_combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][9]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][10]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][11]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][12]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][13]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][14]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][15]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][16]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][17]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][18]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][19]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][20]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][21]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][22]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][23]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][24]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][25]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][26]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][27]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][28]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][29]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][30]~combout ;
wire \reconfigure_ip_inst|wmgmt_readdata[8][31]~combout ;
wire \reconfigure_ip_inst|wmgmt_waitrequest[8]~3_combout ;
wire \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_read~q ;
wire \reconfigure_ip_inst|inst_reconfig_reset_sync|resync_chains[0].sync_r[1]~q ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[0]~0_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[1]~1_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[2]~2_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[3]~3_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[4]~4_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[5]~5_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[6]~6_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[7]~7_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[8]~8_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[9]~9_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[10]~10_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[11]~11_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[12]~12_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[13]~13_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[14]~14_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[15]~15_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_write[0]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_read[0]~0_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[0]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[1]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[2]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[3]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[4]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[5]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[6]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[7]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[8]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[9]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[10]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[11]~0_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[0]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[1]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[2]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[3]~combout ;
wire \reconfigure_ip_inst|basic|a5|pif_interface_sel~q ;
wire \reconfigure_ip_inst|basic|a5|pif_ser_shift_load~q ;
wire \reconfigure_ip_inst|offset.sc_offset|offset_cancellation_av|offset_cancellation_done~1_combout ;
wire \reconfigure_ip_inst|cal_seq|tx_cal_busy~q ;
wire \reconfigure_ip_inst|cal_seq|rx_cal_busy~q ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[16]~16_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[17]~17_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[18]~18_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[19]~19_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[20]~20_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[21]~21_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[22]~22_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[23]~23_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[24]~24_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[25]~25_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[26]~26_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[27]~27_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[28]~28_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[29]~29_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[30]~30_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[31]~31_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_write[1]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_read[1]~1_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[12]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[13]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[14]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[15]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[16]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[17]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[18]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[19]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[20]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[21]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[22]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[23]~1_combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[12]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[13]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[14]~combout ;
wire \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[15]~combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[5]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[4]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[0]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~0_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~2_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~0_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~3_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|lpbk_lock~0_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ;
wire \rtl~3_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ;
wire \rtl~4_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ;
wire \rtl~5_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ;
wire \rtl~6_combout ;
wire \rtl~148_combout ;
wire \rtl~149_combout ;
wire \rtl~14_combout ;
wire \rtl~15_combout ;
wire \rtl~16_combout ;
wire \rtl~17_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ;
wire \rtl~18_combout ;
wire \rtl~19_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~0_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~1_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ;
wire \rtl~20_combout ;
wire \rtl~21_combout ;
wire \rtl~22_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ;
wire \rtl~23_combout ;
wire \rtl~24_combout ;
wire \rtl~26_combout ;
wire \rtl~27_combout ;
wire \rtl~28_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ;
wire \rtl~29_combout ;
wire \rtl~30_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_writedata[4]~q ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ;
wire \rtl~32_combout ;
wire \rtl~33_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|LessThan4~0_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ;
wire \rtl~35_combout ;
wire \rtl~36_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ;
wire \rtl~38_combout ;
wire \rtl~39_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ;
wire \rtl~41_combout ;
wire \rtl~42_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ;
wire \rtl~44_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ;
wire \rtl~45_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ;
wire \rtl~46_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ;
wire \rtl~47_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ;
wire \rtl~48_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ;
wire \rtl~49_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ;
wire \rtl~50_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ;
wire \rtl~51_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ;
wire \rtl~52_combout ;
wire \rtl~150_combout ;
wire \rtl~151_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector5~0_combout ;
wire \reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|inst_rmw_sm|result_data[0]~0_combout ;
wire \rtl~152_combout ;
wire \rtl~153_combout ;
wire \rtl~154_combout ;
wire \rtl~155_combout ;
wire \rtl~156_combout ;
wire \rtl~81_combout ;
wire \rtl~157_combout ;
wire \rtl~158_combout ;
wire \rtl~159_combout ;
wire \rtl~160_combout ;
wire \rtl~161_combout ;
wire \~GND~combout ;
wire \reconfig_from_xcvr[20]~input_o ;
wire \reconfig_from_xcvr[21]~input_o ;
wire \reconfig_from_xcvr[22]~input_o ;
wire \reconfig_from_xcvr[23]~input_o ;
wire \reconfig_from_xcvr[28]~input_o ;
wire \reconfig_from_xcvr[29]~input_o ;
wire \reconfig_from_xcvr[30]~input_o ;
wire \reconfig_from_xcvr[31]~input_o ;
wire \reconfig_from_xcvr[36]~input_o ;
wire \reconfig_from_xcvr[37]~input_o ;
wire \reconfig_from_xcvr[38]~input_o ;
wire \reconfig_from_xcvr[39]~input_o ;
wire \reconfig_from_xcvr[40]~input_o ;
wire \reconfig_from_xcvr[41]~input_o ;
wire \reconfig_from_xcvr[42]~input_o ;
wire \reconfig_from_xcvr[43]~input_o ;
wire \reconfig_from_xcvr[44]~input_o ;
wire \reconfig_from_xcvr[45]~input_o ;
wire \reconfig_from_xcvr[66]~input_o ;
wire \reconfig_from_xcvr[67]~input_o ;
wire \reconfig_from_xcvr[68]~input_o ;
wire \reconfig_from_xcvr[69]~input_o ;
wire \reconfig_from_xcvr[74]~input_o ;
wire \reconfig_from_xcvr[75]~input_o ;
wire \reconfig_from_xcvr[76]~input_o ;
wire \reconfig_from_xcvr[77]~input_o ;
wire \reconfig_from_xcvr[82]~input_o ;
wire \reconfig_from_xcvr[83]~input_o ;
wire \reconfig_from_xcvr[84]~input_o ;
wire \reconfig_from_xcvr[85]~input_o ;
wire \reconfig_from_xcvr[86]~input_o ;
wire \reconfig_from_xcvr[87]~input_o ;
wire \reconfig_from_xcvr[88]~input_o ;
wire \reconfig_from_xcvr[89]~input_o ;
wire \reconfig_from_xcvr[90]~input_o ;
wire \reconfig_from_xcvr[91]~input_o ;
wire \reconfig_mgmt_address[3]~input_o ;
wire \reconfig_mgmt_address[4]~input_o ;
wire \reconfig_mgmt_address[5]~input_o ;
wire \reconfig_mgmt_address[6]~input_o ;
wire \reconfig_mgmt_address[1]~input_o ;
wire \reconfig_mgmt_address[0]~input_o ;
wire \reconfig_mgmt_address[2]~input_o ;
wire \reconfig_mgmt_write~input_o ;
wire \reconfig_mgmt_read~input_o ;
wire \reconfig_mgmt_writedata[0]~input_o ;
wire \reconfig_mgmt_writedata[1]~input_o ;
wire \reconfig_mgmt_writedata[2]~input_o ;
wire \reconfig_mgmt_writedata[3]~input_o ;
wire \reconfig_mif_waitrequest~input_o ;
wire \reconfig_mgmt_writedata[16]~input_o ;
wire \reconfig_from_xcvr[0]~input_o ;
wire \reconfig_from_xcvr[46]~input_o ;
wire \reconfig_mgmt_writedata[17]~input_o ;
wire \reconfig_from_xcvr[1]~input_o ;
wire \reconfig_from_xcvr[47]~input_o ;
wire \reconfig_mgmt_writedata[18]~input_o ;
wire \reconfig_from_xcvr[2]~input_o ;
wire \reconfig_from_xcvr[48]~input_o ;
wire \reconfig_mgmt_writedata[19]~input_o ;
wire \reconfig_from_xcvr[3]~input_o ;
wire \reconfig_from_xcvr[49]~input_o ;
wire \reconfig_mgmt_writedata[20]~input_o ;
wire \reconfig_mgmt_writedata[4]~input_o ;
wire \reconfig_from_xcvr[4]~input_o ;
wire \reconfig_from_xcvr[50]~input_o ;
wire \reconfig_mgmt_writedata[21]~input_o ;
wire \reconfig_mgmt_writedata[5]~input_o ;
wire \reconfig_from_xcvr[5]~input_o ;
wire \reconfig_from_xcvr[51]~input_o ;
wire \reconfig_mgmt_writedata[22]~input_o ;
wire \reconfig_mgmt_writedata[6]~input_o ;
wire \reconfig_from_xcvr[6]~input_o ;
wire \reconfig_from_xcvr[52]~input_o ;
wire \reconfig_mgmt_writedata[23]~input_o ;
wire \reconfig_mgmt_writedata[7]~input_o ;
wire \reconfig_from_xcvr[7]~input_o ;
wire \reconfig_from_xcvr[53]~input_o ;
wire \reconfig_mgmt_writedata[24]~input_o ;
wire \reconfig_mgmt_writedata[8]~input_o ;
wire \reconfig_from_xcvr[8]~input_o ;
wire \reconfig_from_xcvr[54]~input_o ;
wire \reconfig_mgmt_writedata[25]~input_o ;
wire \reconfig_mgmt_writedata[9]~input_o ;
wire \reconfig_from_xcvr[9]~input_o ;
wire \reconfig_from_xcvr[55]~input_o ;
wire \reconfig_mgmt_writedata[26]~input_o ;
wire \reconfig_mgmt_writedata[10]~input_o ;
wire \reconfig_from_xcvr[10]~input_o ;
wire \reconfig_from_xcvr[56]~input_o ;
wire \reconfig_mgmt_writedata[27]~input_o ;
wire \reconfig_mgmt_writedata[11]~input_o ;
wire \reconfig_from_xcvr[11]~input_o ;
wire \reconfig_from_xcvr[57]~input_o ;
wire \reconfig_mgmt_writedata[28]~input_o ;
wire \reconfig_mgmt_writedata[12]~input_o ;
wire \reconfig_from_xcvr[12]~input_o ;
wire \reconfig_from_xcvr[58]~input_o ;
wire \reconfig_mgmt_writedata[29]~input_o ;
wire \reconfig_mgmt_writedata[13]~input_o ;
wire \reconfig_from_xcvr[13]~input_o ;
wire \reconfig_from_xcvr[59]~input_o ;
wire \reconfig_mgmt_writedata[30]~input_o ;
wire \reconfig_mgmt_writedata[14]~input_o ;
wire \reconfig_from_xcvr[14]~input_o ;
wire \reconfig_from_xcvr[60]~input_o ;
wire \reconfig_mgmt_writedata[31]~input_o ;
wire \reconfig_mgmt_writedata[15]~input_o ;
wire \reconfig_from_xcvr[15]~input_o ;
wire \reconfig_from_xcvr[61]~input_o ;
wire \reconfig_mif_readdata[15]~input_o ;
wire \reconfig_mif_readdata[14]~input_o ;
wire \reconfig_mif_readdata[13]~input_o ;
wire \reconfig_mif_readdata[12]~input_o ;
wire \reconfig_mif_readdata[11]~input_o ;
wire \reconfig_mif_readdata[1]~input_o ;
wire \reconfig_mif_readdata[0]~input_o ;
wire \reconfig_mif_readdata[4]~input_o ;
wire \reconfig_mif_readdata[3]~input_o ;
wire \reconfig_mif_readdata[2]~input_o ;
wire \mgmt_rst_reset~input_o ;
wire \reconfig_mif_readdata[7]~input_o ;
wire \reconfig_mif_readdata[5]~input_o ;
wire \reconfig_mif_readdata[6]~input_o ;
wire \reconfig_mif_readdata[8]~input_o ;
wire \reconfig_mif_readdata[9]~input_o ;
wire \reconfig_mif_readdata[10]~input_o ;
wire \reconfig_from_xcvr[24]~input_o ;
wire \reconfig_from_xcvr[70]~input_o ;
wire \reconfig_from_xcvr[16]~input_o ;
wire \reconfig_from_xcvr[62]~input_o ;
wire \reconfig_from_xcvr[32]~input_o ;
wire \reconfig_from_xcvr[78]~input_o ;
wire \reconfig_from_xcvr[25]~input_o ;
wire \reconfig_from_xcvr[71]~input_o ;
wire \reconfig_from_xcvr[17]~input_o ;
wire \reconfig_from_xcvr[63]~input_o ;
wire \reconfig_from_xcvr[33]~input_o ;
wire \reconfig_from_xcvr[79]~input_o ;
wire \reconfig_from_xcvr[26]~input_o ;
wire \reconfig_from_xcvr[72]~input_o ;
wire \reconfig_from_xcvr[18]~input_o ;
wire \reconfig_from_xcvr[64]~input_o ;
wire \reconfig_from_xcvr[34]~input_o ;
wire \reconfig_from_xcvr[80]~input_o ;
wire \reconfig_from_xcvr[27]~input_o ;
wire \reconfig_from_xcvr[73]~input_o ;
wire \reconfig_from_xcvr[19]~input_o ;
wire \reconfig_from_xcvr[65]~input_o ;
wire \reconfig_from_xcvr[35]~input_o ;
wire \reconfig_from_xcvr[81]~input_o ;
wire \mgmt_clk_clk~input_o ;


RECONFIGURE_IP_alt_xcvr_reconfig reconfigure_ip_inst(
	.stream_address_0(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[0]~q ),
	.stream_address_1(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[1]~q ),
	.stream_address_2(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[2]~q ),
	.stream_address_3(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[3]~q ),
	.stream_address_4(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[4]~q ),
	.stream_address_5(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[5]~q ),
	.stream_address_6(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[6]~q ),
	.stream_address_7(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[7]~q ),
	.stream_address_8(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[8]~q ),
	.stream_address_9(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[9]~q ),
	.stream_address_10(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[10]~q ),
	.stream_address_11(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[11]~q ),
	.stream_address_12(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[12]~q ),
	.stream_address_13(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[13]~q ),
	.stream_address_14(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[14]~q ),
	.stream_address_15(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[15]~q ),
	.stream_address_16(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[16]~q ),
	.stream_address_17(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[17]~q ),
	.stream_address_18(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[18]~q ),
	.stream_address_19(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[19]~q ),
	.stream_address_20(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[20]~q ),
	.stream_address_21(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[21]~q ),
	.stream_address_22(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[22]~q ),
	.stream_address_23(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[23]~q ),
	.stream_address_24(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[24]~q ),
	.stream_address_25(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[25]~q ),
	.stream_address_26(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[26]~q ),
	.stream_address_27(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[27]~q ),
	.stream_address_28(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[28]~q ),
	.stream_address_29(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[29]~q ),
	.stream_address_30(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[30]~q ),
	.stream_address_31(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[31]~q ),
	.rtl(\rtl~162_combout ),
	.reconfig_busy(\reconfigure_ip_inst|cal_seq|reconfig_busy~q ),
	.wmgmt_readdata_0_8(\reconfigure_ip_inst|wmgmt_readdata[8][0]~combout ),
	.wmgmt_readdata_1_8(\reconfigure_ip_inst|wmgmt_readdata[8][1]~combout ),
	.wmgmt_readdata_2_8(\reconfigure_ip_inst|wmgmt_readdata[8][2]~combout ),
	.wmgmt_readdata_3_8(\reconfigure_ip_inst|wmgmt_readdata[8][3]~combout ),
	.wmgmt_readdata_4_8(\reconfigure_ip_inst|wmgmt_readdata[8][4]~combout ),
	.wmgmt_readdata_5_8(\reconfigure_ip_inst|wmgmt_readdata[8][5]~combout ),
	.wmgmt_readdata_6_8(\reconfigure_ip_inst|wmgmt_readdata[8][6]~combout ),
	.wmgmt_readdata_7_8(\reconfigure_ip_inst|wmgmt_readdata[8][7]~combout ),
	.reconfig_mgmt_readdata_8(\reconfigure_ip_inst|reconfig_mgmt_readdata[8]~3_combout ),
	.wmgmt_readdata_9_8(\reconfigure_ip_inst|wmgmt_readdata[8][9]~combout ),
	.wmgmt_readdata_10_8(\reconfigure_ip_inst|wmgmt_readdata[8][10]~combout ),
	.wmgmt_readdata_11_8(\reconfigure_ip_inst|wmgmt_readdata[8][11]~combout ),
	.wmgmt_readdata_12_8(\reconfigure_ip_inst|wmgmt_readdata[8][12]~combout ),
	.wmgmt_readdata_13_8(\reconfigure_ip_inst|wmgmt_readdata[8][13]~combout ),
	.wmgmt_readdata_14_8(\reconfigure_ip_inst|wmgmt_readdata[8][14]~combout ),
	.wmgmt_readdata_15_8(\reconfigure_ip_inst|wmgmt_readdata[8][15]~combout ),
	.wmgmt_readdata_16_8(\reconfigure_ip_inst|wmgmt_readdata[8][16]~combout ),
	.wmgmt_readdata_17_8(\reconfigure_ip_inst|wmgmt_readdata[8][17]~combout ),
	.wmgmt_readdata_18_8(\reconfigure_ip_inst|wmgmt_readdata[8][18]~combout ),
	.wmgmt_readdata_19_8(\reconfigure_ip_inst|wmgmt_readdata[8][19]~combout ),
	.wmgmt_readdata_20_8(\reconfigure_ip_inst|wmgmt_readdata[8][20]~combout ),
	.wmgmt_readdata_21_8(\reconfigure_ip_inst|wmgmt_readdata[8][21]~combout ),
	.wmgmt_readdata_22_8(\reconfigure_ip_inst|wmgmt_readdata[8][22]~combout ),
	.wmgmt_readdata_23_8(\reconfigure_ip_inst|wmgmt_readdata[8][23]~combout ),
	.wmgmt_readdata_24_8(\reconfigure_ip_inst|wmgmt_readdata[8][24]~combout ),
	.wmgmt_readdata_25_8(\reconfigure_ip_inst|wmgmt_readdata[8][25]~combout ),
	.wmgmt_readdata_26_8(\reconfigure_ip_inst|wmgmt_readdata[8][26]~combout ),
	.wmgmt_readdata_27_8(\reconfigure_ip_inst|wmgmt_readdata[8][27]~combout ),
	.wmgmt_readdata_28_8(\reconfigure_ip_inst|wmgmt_readdata[8][28]~combout ),
	.wmgmt_readdata_29_8(\reconfigure_ip_inst|wmgmt_readdata[8][29]~combout ),
	.wmgmt_readdata_30_8(\reconfigure_ip_inst|wmgmt_readdata[8][30]~combout ),
	.wmgmt_readdata_31_8(\reconfigure_ip_inst|wmgmt_readdata[8][31]~combout ),
	.wmgmt_waitrequest_8(\reconfigure_ip_inst|wmgmt_waitrequest[8]~3_combout ),
	.stream_read(\reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_read~q ),
	.resync_chains0sync_r_1(\reconfigure_ip_inst|inst_reconfig_reset_sync|resync_chains[0].sync_r[1]~q ),
	.native_reconfig_writedata_0(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[0]~0_combout ),
	.native_reconfig_writedata_1(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[1]~1_combout ),
	.native_reconfig_writedata_2(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[2]~2_combout ),
	.native_reconfig_writedata_3(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[3]~3_combout ),
	.native_reconfig_writedata_4(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[4]~4_combout ),
	.native_reconfig_writedata_5(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[5]~5_combout ),
	.native_reconfig_writedata_6(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[6]~6_combout ),
	.native_reconfig_writedata_7(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[7]~7_combout ),
	.native_reconfig_writedata_8(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[8]~8_combout ),
	.native_reconfig_writedata_9(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[9]~9_combout ),
	.native_reconfig_writedata_10(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[10]~10_combout ),
	.native_reconfig_writedata_11(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[11]~11_combout ),
	.native_reconfig_writedata_12(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[12]~12_combout ),
	.native_reconfig_writedata_13(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[13]~13_combout ),
	.native_reconfig_writedata_14(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[14]~14_combout ),
	.native_reconfig_writedata_15(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[15]~15_combout ),
	.native_reconfig_write_0(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_write[0]~combout ),
	.native_reconfig_read_0(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_read[0]~0_combout ),
	.native_reconfig_address_0(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[0]~combout ),
	.native_reconfig_address_1(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[1]~combout ),
	.native_reconfig_address_2(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[2]~combout ),
	.native_reconfig_address_3(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[3]~combout ),
	.native_reconfig_address_4(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[4]~combout ),
	.native_reconfig_address_5(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[5]~combout ),
	.native_reconfig_address_6(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[6]~combout ),
	.native_reconfig_address_7(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[7]~combout ),
	.native_reconfig_address_8(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[8]~combout ),
	.native_reconfig_address_9(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[9]~combout ),
	.native_reconfig_address_10(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[10]~combout ),
	.native_reconfig_address_11(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[11]~0_combout ),
	.pif_testbus_sel_0(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[0]~combout ),
	.pif_testbus_sel_1(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[1]~combout ),
	.pif_testbus_sel_2(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[2]~combout ),
	.pif_testbus_sel_3(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[3]~combout ),
	.pif_interface_sel(\reconfigure_ip_inst|basic|a5|pif_interface_sel~q ),
	.pif_ser_shift_load(\reconfigure_ip_inst|basic|a5|pif_ser_shift_load~q ),
	.offset_cancellation_done(\reconfigure_ip_inst|offset.sc_offset|offset_cancellation_av|offset_cancellation_done~1_combout ),
	.tx_cal_busy(\reconfigure_ip_inst|cal_seq|tx_cal_busy~q ),
	.rx_cal_busy(\reconfigure_ip_inst|cal_seq|rx_cal_busy~q ),
	.native_reconfig_writedata_16(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[16]~16_combout ),
	.native_reconfig_writedata_17(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[17]~17_combout ),
	.native_reconfig_writedata_18(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[18]~18_combout ),
	.native_reconfig_writedata_19(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[19]~19_combout ),
	.native_reconfig_writedata_20(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[20]~20_combout ),
	.native_reconfig_writedata_21(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[21]~21_combout ),
	.native_reconfig_writedata_22(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[22]~22_combout ),
	.native_reconfig_writedata_23(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[23]~23_combout ),
	.native_reconfig_writedata_24(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[24]~24_combout ),
	.native_reconfig_writedata_25(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[25]~25_combout ),
	.native_reconfig_writedata_26(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[26]~26_combout ),
	.native_reconfig_writedata_27(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[27]~27_combout ),
	.native_reconfig_writedata_28(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[28]~28_combout ),
	.native_reconfig_writedata_29(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[29]~29_combout ),
	.native_reconfig_writedata_30(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[30]~30_combout ),
	.native_reconfig_writedata_31(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[31]~31_combout ),
	.native_reconfig_write_1(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_write[1]~combout ),
	.native_reconfig_read_1(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_read[1]~1_combout ),
	.native_reconfig_address_12(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[12]~combout ),
	.native_reconfig_address_13(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[13]~combout ),
	.native_reconfig_address_14(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[14]~combout ),
	.native_reconfig_address_15(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[15]~combout ),
	.native_reconfig_address_16(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[16]~combout ),
	.native_reconfig_address_17(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[17]~combout ),
	.native_reconfig_address_18(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[18]~combout ),
	.native_reconfig_address_19(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[19]~combout ),
	.native_reconfig_address_20(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[20]~combout ),
	.native_reconfig_address_21(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[21]~combout ),
	.native_reconfig_address_22(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[22]~combout ),
	.native_reconfig_address_23(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[23]~1_combout ),
	.pif_testbus_sel_12(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[12]~combout ),
	.pif_testbus_sel_13(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[13]~combout ),
	.pif_testbus_sel_14(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[14]~combout ),
	.pif_testbus_sel_15(\reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[15]~combout ),
	.uif_addr_offset_5(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[5]~q ),
	.uif_addr_offset_4(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[4]~q ),
	.uif_addr_offset_0(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[0]~q ),
	.Decoder3(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~0_combout ),
	.readdata_for_user_2(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ),
	.readdata_for_user_0(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q ),
	.readdata_for_user_3(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ),
	.readdata_for_user_1(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ),
	.Decoder31(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~2_combout ),
	.Selector2(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~0_combout ),
	.Selector21(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.Decoder32(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~3_combout ),
	.lpbk_lock(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|lpbk_lock~0_combout ),
	.analog_offset_0(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.readdata_for_user_10(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ),
	.readdata_for_user_8(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ),
	.readdata_for_user_11(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ),
	.readdata_for_user_9(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ),
	.rtl1(\rtl~4_combout ),
	.readdata_for_user_6(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ),
	.readdata_for_user_4(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ),
	.readdata_for_user_7(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ),
	.readdata_for_user_5(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ),
	.readdata_for_user_14(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ),
	.readdata_for_user_12(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ),
	.readdata_for_user_15(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ),
	.readdata_for_user_13(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ),
	.rtl2(\rtl~6_combout ),
	.rtl3(\rtl~148_combout ),
	.rtl4(\rtl~149_combout ),
	.rtl5(\rtl~14_combout ),
	.rtl6(\rtl~16_combout ),
	.readdata_for_user_16(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.rtl7(\rtl~18_combout ),
	.rtl8(\rtl~19_combout ),
	.WideOr4(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~0_combout ),
	.WideOr41(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ),
	.analog_length(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.analog_length1(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~1_combout ),
	.analog_length2(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.rtl9(\rtl~21_combout ),
	.readdata_for_user_17(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.rtl10(\rtl~23_combout ),
	.rtl11(\rtl~24_combout ),
	.rtl12(\rtl~27_combout ),
	.readdata_for_user_18(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.rtl13(\rtl~29_combout ),
	.rtl14(\rtl~30_combout ),
	.uif_writedata_4(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_writedata[4]~q ),
	.readdata_for_user_19(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.rtl15(\rtl~32_combout ),
	.rtl16(\rtl~33_combout ),
	.LessThan4(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|LessThan4~0_combout ),
	.readdata_for_user_20(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.rtl17(\rtl~35_combout ),
	.rtl18(\rtl~36_combout ),
	.readdata_for_user_21(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.rtl19(\rtl~38_combout ),
	.rtl20(\rtl~39_combout ),
	.readdata_for_user_22(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.rtl21(\rtl~41_combout ),
	.rtl22(\rtl~42_combout ),
	.readdata_for_user_23(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.rtl23(\rtl~44_combout ),
	.readdata_for_user_24(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.rtl24(\rtl~45_combout ),
	.readdata_for_user_25(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ),
	.rtl25(\rtl~46_combout ),
	.readdata_for_user_26(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ),
	.rtl26(\rtl~47_combout ),
	.readdata_for_user_27(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ),
	.rtl27(\rtl~48_combout ),
	.readdata_for_user_28(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ),
	.rtl28(\rtl~49_combout ),
	.readdata_for_user_29(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ),
	.rtl29(\rtl~50_combout ),
	.readdata_for_user_30(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ),
	.rtl30(\rtl~51_combout ),
	.readdata_for_user_31(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ),
	.rtl31(\rtl~52_combout ),
	.rtl32(\rtl~150_combout ),
	.rtl33(\rtl~151_combout ),
	.Selector5(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector5~0_combout ),
	.result_data_0(\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|inst_rmw_sm|result_data[0]~0_combout ),
	.rtl34(\rtl~153_combout ),
	.rtl35(\rtl~154_combout ),
	.rtl36(\rtl~155_combout ),
	.rtl37(\rtl~156_combout ),
	.rtl38(\rtl~81_combout ),
	.rtl39(\rtl~157_combout ),
	.rtl40(\rtl~158_combout ),
	.rtl41(\rtl~159_combout ),
	.rtl42(\rtl~160_combout ),
	.rtl43(\rtl~161_combout ),
	.GND_port(\~GND~combout ),
	.reconfig_mgmt_address_3(\reconfig_mgmt_address[3]~input_o ),
	.reconfig_mgmt_address_4(\reconfig_mgmt_address[4]~input_o ),
	.reconfig_mgmt_address_5(\reconfig_mgmt_address[5]~input_o ),
	.reconfig_mgmt_address_6(\reconfig_mgmt_address[6]~input_o ),
	.reconfig_mgmt_address_1(\reconfig_mgmt_address[1]~input_o ),
	.reconfig_mgmt_address_0(\reconfig_mgmt_address[0]~input_o ),
	.reconfig_mgmt_address_2(\reconfig_mgmt_address[2]~input_o ),
	.reconfig_mgmt_write(\reconfig_mgmt_write~input_o ),
	.reconfig_mgmt_read(\reconfig_mgmt_read~input_o ),
	.mgmt_clk_clk(\mgmt_clk_clk~input_o ),
	.reconfig_mgmt_writedata_0(\reconfig_mgmt_writedata[0]~input_o ),
	.reconfig_mgmt_writedata_1(\reconfig_mgmt_writedata[1]~input_o ),
	.reconfig_mgmt_writedata_2(\reconfig_mgmt_writedata[2]~input_o ),
	.reconfig_mgmt_writedata_3(\reconfig_mgmt_writedata[3]~input_o ),
	.reconfig_mif_waitrequest(\reconfig_mif_waitrequest~input_o ),
	.reconfig_mgmt_writedata_16(\reconfig_mgmt_writedata[16]~input_o ),
	.reconfig_from_xcvr_0(\reconfig_from_xcvr[0]~input_o ),
	.reconfig_from_xcvr_46(\reconfig_from_xcvr[46]~input_o ),
	.reconfig_mgmt_writedata_17(\reconfig_mgmt_writedata[17]~input_o ),
	.reconfig_from_xcvr_1(\reconfig_from_xcvr[1]~input_o ),
	.reconfig_from_xcvr_47(\reconfig_from_xcvr[47]~input_o ),
	.reconfig_mgmt_writedata_18(\reconfig_mgmt_writedata[18]~input_o ),
	.reconfig_from_xcvr_2(\reconfig_from_xcvr[2]~input_o ),
	.reconfig_from_xcvr_48(\reconfig_from_xcvr[48]~input_o ),
	.reconfig_mgmt_writedata_19(\reconfig_mgmt_writedata[19]~input_o ),
	.reconfig_from_xcvr_3(\reconfig_from_xcvr[3]~input_o ),
	.reconfig_from_xcvr_49(\reconfig_from_xcvr[49]~input_o ),
	.reconfig_mgmt_writedata_20(\reconfig_mgmt_writedata[20]~input_o ),
	.reconfig_mgmt_writedata_4(\reconfig_mgmt_writedata[4]~input_o ),
	.reconfig_from_xcvr_4(\reconfig_from_xcvr[4]~input_o ),
	.reconfig_from_xcvr_50(\reconfig_from_xcvr[50]~input_o ),
	.reconfig_mgmt_writedata_21(\reconfig_mgmt_writedata[21]~input_o ),
	.reconfig_mgmt_writedata_5(\reconfig_mgmt_writedata[5]~input_o ),
	.reconfig_from_xcvr_5(\reconfig_from_xcvr[5]~input_o ),
	.reconfig_from_xcvr_51(\reconfig_from_xcvr[51]~input_o ),
	.reconfig_mgmt_writedata_22(\reconfig_mgmt_writedata[22]~input_o ),
	.reconfig_mgmt_writedata_6(\reconfig_mgmt_writedata[6]~input_o ),
	.reconfig_from_xcvr_6(\reconfig_from_xcvr[6]~input_o ),
	.reconfig_from_xcvr_52(\reconfig_from_xcvr[52]~input_o ),
	.reconfig_mgmt_writedata_23(\reconfig_mgmt_writedata[23]~input_o ),
	.reconfig_mgmt_writedata_7(\reconfig_mgmt_writedata[7]~input_o ),
	.reconfig_from_xcvr_7(\reconfig_from_xcvr[7]~input_o ),
	.reconfig_from_xcvr_53(\reconfig_from_xcvr[53]~input_o ),
	.reconfig_mgmt_writedata_24(\reconfig_mgmt_writedata[24]~input_o ),
	.reconfig_mgmt_writedata_8(\reconfig_mgmt_writedata[8]~input_o ),
	.reconfig_from_xcvr_8(\reconfig_from_xcvr[8]~input_o ),
	.reconfig_from_xcvr_54(\reconfig_from_xcvr[54]~input_o ),
	.reconfig_mgmt_writedata_25(\reconfig_mgmt_writedata[25]~input_o ),
	.reconfig_mgmt_writedata_9(\reconfig_mgmt_writedata[9]~input_o ),
	.reconfig_from_xcvr_9(\reconfig_from_xcvr[9]~input_o ),
	.reconfig_from_xcvr_55(\reconfig_from_xcvr[55]~input_o ),
	.reconfig_mgmt_writedata_26(\reconfig_mgmt_writedata[26]~input_o ),
	.reconfig_mgmt_writedata_10(\reconfig_mgmt_writedata[10]~input_o ),
	.reconfig_from_xcvr_10(\reconfig_from_xcvr[10]~input_o ),
	.reconfig_from_xcvr_56(\reconfig_from_xcvr[56]~input_o ),
	.reconfig_mgmt_writedata_27(\reconfig_mgmt_writedata[27]~input_o ),
	.reconfig_mgmt_writedata_11(\reconfig_mgmt_writedata[11]~input_o ),
	.reconfig_from_xcvr_11(\reconfig_from_xcvr[11]~input_o ),
	.reconfig_from_xcvr_57(\reconfig_from_xcvr[57]~input_o ),
	.reconfig_mgmt_writedata_28(\reconfig_mgmt_writedata[28]~input_o ),
	.reconfig_mgmt_writedata_12(\reconfig_mgmt_writedata[12]~input_o ),
	.reconfig_from_xcvr_12(\reconfig_from_xcvr[12]~input_o ),
	.reconfig_from_xcvr_58(\reconfig_from_xcvr[58]~input_o ),
	.reconfig_mgmt_writedata_29(\reconfig_mgmt_writedata[29]~input_o ),
	.reconfig_mgmt_writedata_13(\reconfig_mgmt_writedata[13]~input_o ),
	.reconfig_from_xcvr_13(\reconfig_from_xcvr[13]~input_o ),
	.reconfig_from_xcvr_59(\reconfig_from_xcvr[59]~input_o ),
	.reconfig_mgmt_writedata_30(\reconfig_mgmt_writedata[30]~input_o ),
	.reconfig_mgmt_writedata_14(\reconfig_mgmt_writedata[14]~input_o ),
	.reconfig_from_xcvr_14(\reconfig_from_xcvr[14]~input_o ),
	.reconfig_from_xcvr_60(\reconfig_from_xcvr[60]~input_o ),
	.reconfig_mgmt_writedata_31(\reconfig_mgmt_writedata[31]~input_o ),
	.reconfig_mgmt_writedata_15(\reconfig_mgmt_writedata[15]~input_o ),
	.reconfig_from_xcvr_15(\reconfig_from_xcvr[15]~input_o ),
	.reconfig_from_xcvr_61(\reconfig_from_xcvr[61]~input_o ),
	.reconfig_mif_readdata_15(\reconfig_mif_readdata[15]~input_o ),
	.reconfig_mif_readdata_14(\reconfig_mif_readdata[14]~input_o ),
	.reconfig_mif_readdata_13(\reconfig_mif_readdata[13]~input_o ),
	.reconfig_mif_readdata_12(\reconfig_mif_readdata[12]~input_o ),
	.reconfig_mif_readdata_11(\reconfig_mif_readdata[11]~input_o ),
	.reconfig_mif_readdata_1(\reconfig_mif_readdata[1]~input_o ),
	.reconfig_mif_readdata_0(\reconfig_mif_readdata[0]~input_o ),
	.reconfig_mif_readdata_4(\reconfig_mif_readdata[4]~input_o ),
	.reconfig_mif_readdata_3(\reconfig_mif_readdata[3]~input_o ),
	.reconfig_mif_readdata_2(\reconfig_mif_readdata[2]~input_o ),
	.mgmt_rst_reset(\mgmt_rst_reset~input_o ),
	.reconfig_mif_readdata_7(\reconfig_mif_readdata[7]~input_o ),
	.reconfig_mif_readdata_5(\reconfig_mif_readdata[5]~input_o ),
	.reconfig_mif_readdata_6(\reconfig_mif_readdata[6]~input_o ),
	.reconfig_mif_readdata_8(\reconfig_mif_readdata[8]~input_o ),
	.reconfig_mif_readdata_9(\reconfig_mif_readdata[9]~input_o ),
	.reconfig_mif_readdata_10(\reconfig_mif_readdata[10]~input_o ),
	.reconfig_from_xcvr_24(\reconfig_from_xcvr[24]~input_o ),
	.reconfig_from_xcvr_70(\reconfig_from_xcvr[70]~input_o ),
	.reconfig_from_xcvr_16(\reconfig_from_xcvr[16]~input_o ),
	.reconfig_from_xcvr_62(\reconfig_from_xcvr[62]~input_o ),
	.reconfig_from_xcvr_32(\reconfig_from_xcvr[32]~input_o ),
	.reconfig_from_xcvr_78(\reconfig_from_xcvr[78]~input_o ),
	.reconfig_from_xcvr_25(\reconfig_from_xcvr[25]~input_o ),
	.reconfig_from_xcvr_71(\reconfig_from_xcvr[71]~input_o ),
	.reconfig_from_xcvr_17(\reconfig_from_xcvr[17]~input_o ),
	.reconfig_from_xcvr_63(\reconfig_from_xcvr[63]~input_o ),
	.reconfig_from_xcvr_33(\reconfig_from_xcvr[33]~input_o ),
	.reconfig_from_xcvr_79(\reconfig_from_xcvr[79]~input_o ),
	.reconfig_from_xcvr_26(\reconfig_from_xcvr[26]~input_o ),
	.reconfig_from_xcvr_72(\reconfig_from_xcvr[72]~input_o ),
	.reconfig_from_xcvr_18(\reconfig_from_xcvr[18]~input_o ),
	.reconfig_from_xcvr_64(\reconfig_from_xcvr[64]~input_o ),
	.reconfig_from_xcvr_34(\reconfig_from_xcvr[34]~input_o ),
	.reconfig_from_xcvr_80(\reconfig_from_xcvr[80]~input_o ),
	.reconfig_from_xcvr_27(\reconfig_from_xcvr[27]~input_o ),
	.reconfig_from_xcvr_73(\reconfig_from_xcvr[73]~input_o ),
	.reconfig_from_xcvr_19(\reconfig_from_xcvr[19]~input_o ),
	.reconfig_from_xcvr_65(\reconfig_from_xcvr[65]~input_o ),
	.reconfig_from_xcvr_35(\reconfig_from_xcvr[35]~input_o ),
	.reconfig_from_xcvr_81(\reconfig_from_xcvr[81]~input_o ));

cyclonev_lcell_comb \rtl~162 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[5]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.datac(!\rtl~152_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector5~0_combout ),
	.datag(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~2_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~162_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~162 .extended_lut = "on";
defparam \rtl~162 .lut_mask = 64'h00000F0F020A0F0F;
defparam \rtl~162 .shared_arith = "off";

cyclonev_lcell_comb \rtl~3 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~3 .extended_lut = "off";
defparam \rtl~3 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~3 .shared_arith = "off";

cyclonev_lcell_comb \rtl~4 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~4 .extended_lut = "off";
defparam \rtl~4 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~4 .shared_arith = "off";

cyclonev_lcell_comb \rtl~5 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~5 .extended_lut = "off";
defparam \rtl~5 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~5 .shared_arith = "off";

cyclonev_lcell_comb \rtl~6 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~6 .extended_lut = "off";
defparam \rtl~6 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~6 .shared_arith = "off";

cyclonev_lcell_comb \rtl~148 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[5]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[4]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[0]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~0_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|lpbk_lock~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~148_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~148 .extended_lut = "off";
defparam \rtl~148 .lut_mask = 64'h0004004600040046;
defparam \rtl~148 .shared_arith = "off";

cyclonev_lcell_comb \rtl~149 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[5]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[4]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_addr_offset[0]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~0_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|lpbk_lock~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~149_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~149 .extended_lut = "off";
defparam \rtl~149 .lut_mask = 64'h0084008200840082;
defparam \rtl~149 .shared_arith = "off";

cyclonev_lcell_comb \rtl~14 (
	.dataa(!\rtl~3_combout ),
	.datab(!\rtl~4_combout ),
	.datac(!\rtl~5_combout ),
	.datad(!\rtl~6_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~14 .extended_lut = "off";
defparam \rtl~14 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~14 .shared_arith = "off";

cyclonev_lcell_comb \rtl~15 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~15 .extended_lut = "off";
defparam \rtl~15 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~15 .shared_arith = "off";

cyclonev_lcell_comb \rtl~16 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~16 .extended_lut = "off";
defparam \rtl~16 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~16 .shared_arith = "off";

cyclonev_lcell_comb \rtl~17 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~17 .extended_lut = "off";
defparam \rtl~17 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~17 .shared_arith = "off";

cyclonev_lcell_comb \rtl~18 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~18 .extended_lut = "off";
defparam \rtl~18 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~18 .shared_arith = "off";

cyclonev_lcell_comb \rtl~19 (
	.dataa(!\rtl~15_combout ),
	.datab(!\rtl~16_combout ),
	.datac(!\rtl~17_combout ),
	.datad(!\rtl~18_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~19 .extended_lut = "off";
defparam \rtl~19 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~19 .shared_arith = "off";

cyclonev_lcell_comb \rtl~20 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~20 .extended_lut = "off";
defparam \rtl~20 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~20 .shared_arith = "off";

cyclonev_lcell_comb \rtl~21 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~21 .extended_lut = "off";
defparam \rtl~21 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~21 .shared_arith = "off";

cyclonev_lcell_comb \rtl~22 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~22 .extended_lut = "off";
defparam \rtl~22 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~22 .shared_arith = "off";

cyclonev_lcell_comb \rtl~23 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~23 .extended_lut = "off";
defparam \rtl~23 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~23 .shared_arith = "off";

cyclonev_lcell_comb \rtl~24 (
	.dataa(!\rtl~20_combout ),
	.datab(!\rtl~21_combout ),
	.datac(!\rtl~22_combout ),
	.datad(!\rtl~23_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~24 .extended_lut = "off";
defparam \rtl~24 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~24 .shared_arith = "off";

cyclonev_lcell_comb \rtl~26 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~26 .extended_lut = "off";
defparam \rtl~26 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~26 .shared_arith = "off";

cyclonev_lcell_comb \rtl~27 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~27 .extended_lut = "off";
defparam \rtl~27 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~27 .shared_arith = "off";

cyclonev_lcell_comb \rtl~28 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~28 .extended_lut = "off";
defparam \rtl~28 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~28 .shared_arith = "off";

cyclonev_lcell_comb \rtl~29 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~29 .extended_lut = "off";
defparam \rtl~29 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~29 .shared_arith = "off";

cyclonev_lcell_comb \rtl~30 (
	.dataa(!\rtl~26_combout ),
	.datab(!\rtl~27_combout ),
	.datac(!\rtl~28_combout ),
	.datad(!\rtl~29_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~30 .extended_lut = "off";
defparam \rtl~30 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~30 .shared_arith = "off";

cyclonev_lcell_comb \rtl~32 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~32 .extended_lut = "off";
defparam \rtl~32 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~32 .shared_arith = "off";

cyclonev_lcell_comb \rtl~33 (
	.dataa(!\rtl~5_combout ),
	.datab(!\rtl~6_combout ),
	.datac(!\rtl~4_combout ),
	.datad(!\rtl~32_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~33 .extended_lut = "off";
defparam \rtl~33 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~33 .shared_arith = "off";

cyclonev_lcell_comb \rtl~35 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~35 .extended_lut = "off";
defparam \rtl~35 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~35 .shared_arith = "off";

cyclonev_lcell_comb \rtl~36 (
	.dataa(!\rtl~17_combout ),
	.datab(!\rtl~18_combout ),
	.datac(!\rtl~16_combout ),
	.datad(!\rtl~35_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~36 .extended_lut = "off";
defparam \rtl~36 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~36 .shared_arith = "off";

cyclonev_lcell_comb \rtl~38 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~38 .extended_lut = "off";
defparam \rtl~38 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~38 .shared_arith = "off";

cyclonev_lcell_comb \rtl~39 (
	.dataa(!\rtl~22_combout ),
	.datab(!\rtl~23_combout ),
	.datac(!\rtl~21_combout ),
	.datad(!\rtl~38_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~39 .extended_lut = "off";
defparam \rtl~39 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~39 .shared_arith = "off";

cyclonev_lcell_comb \rtl~41 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~41 .extended_lut = "off";
defparam \rtl~41 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~41 .shared_arith = "off";

cyclonev_lcell_comb \rtl~42 (
	.dataa(!\rtl~28_combout ),
	.datab(!\rtl~29_combout ),
	.datac(!\rtl~27_combout ),
	.datad(!\rtl~41_combout ),
	.datae(!\rtl~148_combout ),
	.dataf(!\rtl~149_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~42 .extended_lut = "off";
defparam \rtl~42 .lut_mask = 64'h555533330F0F00FF;
defparam \rtl~42 .shared_arith = "off";

cyclonev_lcell_comb \rtl~44 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~44 .extended_lut = "off";
defparam \rtl~44 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~44 .shared_arith = "off";

cyclonev_lcell_comb \rtl~45 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~45 .extended_lut = "off";
defparam \rtl~45 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~45 .shared_arith = "off";

cyclonev_lcell_comb \rtl~46 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~46 .extended_lut = "off";
defparam \rtl~46 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~46 .shared_arith = "off";

cyclonev_lcell_comb \rtl~47 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~47 .extended_lut = "off";
defparam \rtl~47 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~47 .shared_arith = "off";

cyclonev_lcell_comb \rtl~48 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~48 .extended_lut = "off";
defparam \rtl~48 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~48 .shared_arith = "off";

cyclonev_lcell_comb \rtl~49 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~49 .extended_lut = "off";
defparam \rtl~49 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~49 .shared_arith = "off";

cyclonev_lcell_comb \rtl~50 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~50 .extended_lut = "off";
defparam \rtl~50 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~50 .shared_arith = "off";

cyclonev_lcell_comb \rtl~51 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~51 .extended_lut = "off";
defparam \rtl~51 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~51 .shared_arith = "off";

cyclonev_lcell_comb \rtl~52 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~52 .extended_lut = "off";
defparam \rtl~52 .lut_mask = 64'h3333555500FF0F0F;
defparam \rtl~52 .shared_arith = "off";

cyclonev_lcell_comb \rtl~150 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~150_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~150 .extended_lut = "off";
defparam \rtl~150 .lut_mask = 64'h084C2A6E084C2A6E;
defparam \rtl~150 .shared_arith = "off";

cyclonev_lcell_comb \rtl~151 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~2_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~3_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|lpbk_lock~0_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~0_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~151_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~151 .extended_lut = "off";
defparam \rtl~151 .lut_mask = 64'h0000CF8A3020FFAA;
defparam \rtl~151 .shared_arith = "off";

cyclonev_lcell_comb \rtl~152 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|inst_rmw_sm|result_data[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~152_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~152 .extended_lut = "off";
defparam \rtl~152 .lut_mask = 64'h007F007F007F007F;
defparam \rtl~152 .shared_arith = "off";

cyclonev_lcell_comb \rtl~153 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~153_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~153 .extended_lut = "off";
defparam \rtl~153 .lut_mask = 64'hE000E000E000E000;
defparam \rtl~153 .shared_arith = "off";

cyclonev_lcell_comb \rtl~154 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datac(!\rtl~152_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~154_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~154 .extended_lut = "off";
defparam \rtl~154 .lut_mask = 64'h0202020202020202;
defparam \rtl~154 .shared_arith = "off";

cyclonev_lcell_comb \rtl~155 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~155_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~155 .extended_lut = "off";
defparam \rtl~155 .lut_mask = 64'h02AA2AAA02AA2AAA;
defparam \rtl~155 .shared_arith = "off";

cyclonev_lcell_comb \rtl~156 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datab(!\rtl~162_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~156_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~156 .extended_lut = "off";
defparam \rtl~156 .lut_mask = 64'h1111111111111111;
defparam \rtl~156 .shared_arith = "off";

cyclonev_lcell_comb \rtl~81 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Decoder3~3_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|lpbk_lock~0_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.dataf(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~81 .extended_lut = "off";
defparam \rtl~81 .lut_mask = 64'hFFEFEF0000000000;
defparam \rtl~81 .shared_arith = "off";

cyclonev_lcell_comb \rtl~157 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~157_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~157 .extended_lut = "off";
defparam \rtl~157 .lut_mask = 64'h0000000200000002;
defparam \rtl~157 .shared_arith = "off";

cyclonev_lcell_comb \rtl~158 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~1_combout ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datae(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~158_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~158 .extended_lut = "off";
defparam \rtl~158 .lut_mask = 64'h0022022200220222;
defparam \rtl~158 .shared_arith = "off";

cyclonev_lcell_comb \rtl~159 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_offset[0]~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_writedata[4]~q ),
	.datad(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|LessThan4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~159_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~159 .extended_lut = "off";
defparam \rtl~159 .lut_mask = 64'h0002000200020002;
defparam \rtl~159 .shared_arith = "off";

cyclonev_lcell_comb \rtl~160 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|Selector2~1_combout ),
	.datab(!\rtl~162_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~160_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~160 .extended_lut = "off";
defparam \rtl~160 .lut_mask = 64'h2222222222222222;
defparam \rtl~160 .shared_arith = "off";

cyclonev_lcell_comb \rtl~161 (
	.dataa(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|WideOr4~0_combout ),
	.datab(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~0_combout ),
	.datac(!\reconfigure_ip_inst|analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|analog_length~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rtl~161_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rtl~161 .extended_lut = "off";
defparam \rtl~161 .lut_mask = 64'h1313131313131313;
defparam \rtl~161 .shared_arith = "off";

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

assign \reconfig_mgmt_address[3]~input_o  = reconfig_mgmt_address[3];

assign \reconfig_mgmt_address[4]~input_o  = reconfig_mgmt_address[4];

assign \reconfig_mgmt_address[5]~input_o  = reconfig_mgmt_address[5];

assign \reconfig_mgmt_address[6]~input_o  = reconfig_mgmt_address[6];

assign \reconfig_mgmt_address[1]~input_o  = reconfig_mgmt_address[1];

assign \reconfig_mgmt_address[0]~input_o  = reconfig_mgmt_address[0];

assign \reconfig_mgmt_address[2]~input_o  = reconfig_mgmt_address[2];

assign \reconfig_mgmt_write~input_o  = reconfig_mgmt_write;

assign \reconfig_mgmt_read~input_o  = reconfig_mgmt_read;

assign \reconfig_mgmt_writedata[0]~input_o  = reconfig_mgmt_writedata[0];

assign \reconfig_mgmt_writedata[1]~input_o  = reconfig_mgmt_writedata[1];

assign \reconfig_mgmt_writedata[2]~input_o  = reconfig_mgmt_writedata[2];

assign \reconfig_mgmt_writedata[3]~input_o  = reconfig_mgmt_writedata[3];

assign \reconfig_mif_waitrequest~input_o  = reconfig_mif_waitrequest;

assign \reconfig_mgmt_writedata[16]~input_o  = reconfig_mgmt_writedata[16];

assign \reconfig_from_xcvr[0]~input_o  = reconfig_from_xcvr[0];

assign \reconfig_from_xcvr[46]~input_o  = reconfig_from_xcvr[46];

assign \reconfig_mgmt_writedata[17]~input_o  = reconfig_mgmt_writedata[17];

assign \reconfig_from_xcvr[1]~input_o  = reconfig_from_xcvr[1];

assign \reconfig_from_xcvr[47]~input_o  = reconfig_from_xcvr[47];

assign \reconfig_mgmt_writedata[18]~input_o  = reconfig_mgmt_writedata[18];

assign \reconfig_from_xcvr[2]~input_o  = reconfig_from_xcvr[2];

assign \reconfig_from_xcvr[48]~input_o  = reconfig_from_xcvr[48];

assign \reconfig_mgmt_writedata[19]~input_o  = reconfig_mgmt_writedata[19];

assign \reconfig_from_xcvr[3]~input_o  = reconfig_from_xcvr[3];

assign \reconfig_from_xcvr[49]~input_o  = reconfig_from_xcvr[49];

assign \reconfig_mgmt_writedata[20]~input_o  = reconfig_mgmt_writedata[20];

assign \reconfig_mgmt_writedata[4]~input_o  = reconfig_mgmt_writedata[4];

assign \reconfig_from_xcvr[4]~input_o  = reconfig_from_xcvr[4];

assign \reconfig_from_xcvr[50]~input_o  = reconfig_from_xcvr[50];

assign \reconfig_mgmt_writedata[21]~input_o  = reconfig_mgmt_writedata[21];

assign \reconfig_mgmt_writedata[5]~input_o  = reconfig_mgmt_writedata[5];

assign \reconfig_from_xcvr[5]~input_o  = reconfig_from_xcvr[5];

assign \reconfig_from_xcvr[51]~input_o  = reconfig_from_xcvr[51];

assign \reconfig_mgmt_writedata[22]~input_o  = reconfig_mgmt_writedata[22];

assign \reconfig_mgmt_writedata[6]~input_o  = reconfig_mgmt_writedata[6];

assign \reconfig_from_xcvr[6]~input_o  = reconfig_from_xcvr[6];

assign \reconfig_from_xcvr[52]~input_o  = reconfig_from_xcvr[52];

assign \reconfig_mgmt_writedata[23]~input_o  = reconfig_mgmt_writedata[23];

assign \reconfig_mgmt_writedata[7]~input_o  = reconfig_mgmt_writedata[7];

assign \reconfig_from_xcvr[7]~input_o  = reconfig_from_xcvr[7];

assign \reconfig_from_xcvr[53]~input_o  = reconfig_from_xcvr[53];

assign \reconfig_mgmt_writedata[24]~input_o  = reconfig_mgmt_writedata[24];

assign \reconfig_mgmt_writedata[8]~input_o  = reconfig_mgmt_writedata[8];

assign \reconfig_from_xcvr[8]~input_o  = reconfig_from_xcvr[8];

assign \reconfig_from_xcvr[54]~input_o  = reconfig_from_xcvr[54];

assign \reconfig_mgmt_writedata[25]~input_o  = reconfig_mgmt_writedata[25];

assign \reconfig_mgmt_writedata[9]~input_o  = reconfig_mgmt_writedata[9];

assign \reconfig_from_xcvr[9]~input_o  = reconfig_from_xcvr[9];

assign \reconfig_from_xcvr[55]~input_o  = reconfig_from_xcvr[55];

assign \reconfig_mgmt_writedata[26]~input_o  = reconfig_mgmt_writedata[26];

assign \reconfig_mgmt_writedata[10]~input_o  = reconfig_mgmt_writedata[10];

assign \reconfig_from_xcvr[10]~input_o  = reconfig_from_xcvr[10];

assign \reconfig_from_xcvr[56]~input_o  = reconfig_from_xcvr[56];

assign \reconfig_mgmt_writedata[27]~input_o  = reconfig_mgmt_writedata[27];

assign \reconfig_mgmt_writedata[11]~input_o  = reconfig_mgmt_writedata[11];

assign \reconfig_from_xcvr[11]~input_o  = reconfig_from_xcvr[11];

assign \reconfig_from_xcvr[57]~input_o  = reconfig_from_xcvr[57];

assign \reconfig_mgmt_writedata[28]~input_o  = reconfig_mgmt_writedata[28];

assign \reconfig_mgmt_writedata[12]~input_o  = reconfig_mgmt_writedata[12];

assign \reconfig_from_xcvr[12]~input_o  = reconfig_from_xcvr[12];

assign \reconfig_from_xcvr[58]~input_o  = reconfig_from_xcvr[58];

assign \reconfig_mgmt_writedata[29]~input_o  = reconfig_mgmt_writedata[29];

assign \reconfig_mgmt_writedata[13]~input_o  = reconfig_mgmt_writedata[13];

assign \reconfig_from_xcvr[13]~input_o  = reconfig_from_xcvr[13];

assign \reconfig_from_xcvr[59]~input_o  = reconfig_from_xcvr[59];

assign \reconfig_mgmt_writedata[30]~input_o  = reconfig_mgmt_writedata[30];

assign \reconfig_mgmt_writedata[14]~input_o  = reconfig_mgmt_writedata[14];

assign \reconfig_from_xcvr[14]~input_o  = reconfig_from_xcvr[14];

assign \reconfig_from_xcvr[60]~input_o  = reconfig_from_xcvr[60];

assign \reconfig_mgmt_writedata[31]~input_o  = reconfig_mgmt_writedata[31];

assign \reconfig_mgmt_writedata[15]~input_o  = reconfig_mgmt_writedata[15];

assign \reconfig_from_xcvr[15]~input_o  = reconfig_from_xcvr[15];

assign \reconfig_from_xcvr[61]~input_o  = reconfig_from_xcvr[61];

assign \reconfig_mif_readdata[15]~input_o  = reconfig_mif_readdata[15];

assign \reconfig_mif_readdata[14]~input_o  = reconfig_mif_readdata[14];

assign \reconfig_mif_readdata[13]~input_o  = reconfig_mif_readdata[13];

assign \reconfig_mif_readdata[12]~input_o  = reconfig_mif_readdata[12];

assign \reconfig_mif_readdata[11]~input_o  = reconfig_mif_readdata[11];

assign \reconfig_mif_readdata[1]~input_o  = reconfig_mif_readdata[1];

assign \reconfig_mif_readdata[0]~input_o  = reconfig_mif_readdata[0];

assign \reconfig_mif_readdata[4]~input_o  = reconfig_mif_readdata[4];

assign \reconfig_mif_readdata[3]~input_o  = reconfig_mif_readdata[3];

assign \reconfig_mif_readdata[2]~input_o  = reconfig_mif_readdata[2];

assign \mgmt_rst_reset~input_o  = mgmt_rst_reset;

assign \reconfig_mif_readdata[7]~input_o  = reconfig_mif_readdata[7];

assign \reconfig_mif_readdata[5]~input_o  = reconfig_mif_readdata[5];

assign \reconfig_mif_readdata[6]~input_o  = reconfig_mif_readdata[6];

assign \reconfig_mif_readdata[8]~input_o  = reconfig_mif_readdata[8];

assign \reconfig_mif_readdata[9]~input_o  = reconfig_mif_readdata[9];

assign \reconfig_mif_readdata[10]~input_o  = reconfig_mif_readdata[10];

assign \reconfig_from_xcvr[24]~input_o  = reconfig_from_xcvr[24];

assign \reconfig_from_xcvr[70]~input_o  = reconfig_from_xcvr[70];

assign \reconfig_from_xcvr[16]~input_o  = reconfig_from_xcvr[16];

assign \reconfig_from_xcvr[62]~input_o  = reconfig_from_xcvr[62];

assign \reconfig_from_xcvr[32]~input_o  = reconfig_from_xcvr[32];

assign \reconfig_from_xcvr[78]~input_o  = reconfig_from_xcvr[78];

assign \reconfig_from_xcvr[25]~input_o  = reconfig_from_xcvr[25];

assign \reconfig_from_xcvr[71]~input_o  = reconfig_from_xcvr[71];

assign \reconfig_from_xcvr[17]~input_o  = reconfig_from_xcvr[17];

assign \reconfig_from_xcvr[63]~input_o  = reconfig_from_xcvr[63];

assign \reconfig_from_xcvr[33]~input_o  = reconfig_from_xcvr[33];

assign \reconfig_from_xcvr[79]~input_o  = reconfig_from_xcvr[79];

assign \reconfig_from_xcvr[26]~input_o  = reconfig_from_xcvr[26];

assign \reconfig_from_xcvr[72]~input_o  = reconfig_from_xcvr[72];

assign \reconfig_from_xcvr[18]~input_o  = reconfig_from_xcvr[18];

assign \reconfig_from_xcvr[64]~input_o  = reconfig_from_xcvr[64];

assign \reconfig_from_xcvr[34]~input_o  = reconfig_from_xcvr[34];

assign \reconfig_from_xcvr[80]~input_o  = reconfig_from_xcvr[80];

assign \reconfig_from_xcvr[27]~input_o  = reconfig_from_xcvr[27];

assign \reconfig_from_xcvr[73]~input_o  = reconfig_from_xcvr[73];

assign \reconfig_from_xcvr[19]~input_o  = reconfig_from_xcvr[19];

assign \reconfig_from_xcvr[65]~input_o  = reconfig_from_xcvr[65];

assign \reconfig_from_xcvr[35]~input_o  = reconfig_from_xcvr[35];

assign \reconfig_from_xcvr[81]~input_o  = reconfig_from_xcvr[81];

assign reconfig_busy = ~ \reconfigure_ip_inst|cal_seq|reconfig_busy~q ;

assign reconfig_mgmt_readdata[0] = \reconfigure_ip_inst|wmgmt_readdata[8][0]~combout ;

assign reconfig_mgmt_readdata[1] = \reconfigure_ip_inst|wmgmt_readdata[8][1]~combout ;

assign reconfig_mgmt_readdata[2] = \reconfigure_ip_inst|wmgmt_readdata[8][2]~combout ;

assign reconfig_mgmt_readdata[3] = \reconfigure_ip_inst|wmgmt_readdata[8][3]~combout ;

assign reconfig_mgmt_readdata[4] = \reconfigure_ip_inst|wmgmt_readdata[8][4]~combout ;

assign reconfig_mgmt_readdata[5] = \reconfigure_ip_inst|wmgmt_readdata[8][5]~combout ;

assign reconfig_mgmt_readdata[6] = \reconfigure_ip_inst|wmgmt_readdata[8][6]~combout ;

assign reconfig_mgmt_readdata[7] = \reconfigure_ip_inst|wmgmt_readdata[8][7]~combout ;

assign reconfig_mgmt_readdata[8] = \reconfigure_ip_inst|reconfig_mgmt_readdata[8]~3_combout ;

assign reconfig_mgmt_readdata[9] = \reconfigure_ip_inst|wmgmt_readdata[8][9]~combout ;

assign reconfig_mgmt_readdata[10] = \reconfigure_ip_inst|wmgmt_readdata[8][10]~combout ;

assign reconfig_mgmt_readdata[11] = \reconfigure_ip_inst|wmgmt_readdata[8][11]~combout ;

assign reconfig_mgmt_readdata[12] = \reconfigure_ip_inst|wmgmt_readdata[8][12]~combout ;

assign reconfig_mgmt_readdata[13] = \reconfigure_ip_inst|wmgmt_readdata[8][13]~combout ;

assign reconfig_mgmt_readdata[14] = \reconfigure_ip_inst|wmgmt_readdata[8][14]~combout ;

assign reconfig_mgmt_readdata[15] = \reconfigure_ip_inst|wmgmt_readdata[8][15]~combout ;

assign reconfig_mgmt_readdata[16] = \reconfigure_ip_inst|wmgmt_readdata[8][16]~combout ;

assign reconfig_mgmt_readdata[17] = \reconfigure_ip_inst|wmgmt_readdata[8][17]~combout ;

assign reconfig_mgmt_readdata[18] = \reconfigure_ip_inst|wmgmt_readdata[8][18]~combout ;

assign reconfig_mgmt_readdata[19] = \reconfigure_ip_inst|wmgmt_readdata[8][19]~combout ;

assign reconfig_mgmt_readdata[20] = \reconfigure_ip_inst|wmgmt_readdata[8][20]~combout ;

assign reconfig_mgmt_readdata[21] = \reconfigure_ip_inst|wmgmt_readdata[8][21]~combout ;

assign reconfig_mgmt_readdata[22] = \reconfigure_ip_inst|wmgmt_readdata[8][22]~combout ;

assign reconfig_mgmt_readdata[23] = \reconfigure_ip_inst|wmgmt_readdata[8][23]~combout ;

assign reconfig_mgmt_readdata[24] = \reconfigure_ip_inst|wmgmt_readdata[8][24]~combout ;

assign reconfig_mgmt_readdata[25] = \reconfigure_ip_inst|wmgmt_readdata[8][25]~combout ;

assign reconfig_mgmt_readdata[26] = \reconfigure_ip_inst|wmgmt_readdata[8][26]~combout ;

assign reconfig_mgmt_readdata[27] = \reconfigure_ip_inst|wmgmt_readdata[8][27]~combout ;

assign reconfig_mgmt_readdata[28] = \reconfigure_ip_inst|wmgmt_readdata[8][28]~combout ;

assign reconfig_mgmt_readdata[29] = \reconfigure_ip_inst|wmgmt_readdata[8][29]~combout ;

assign reconfig_mgmt_readdata[30] = \reconfigure_ip_inst|wmgmt_readdata[8][30]~combout ;

assign reconfig_mgmt_readdata[31] = \reconfigure_ip_inst|wmgmt_readdata[8][31]~combout ;

assign reconfig_mgmt_waitrequest = \reconfigure_ip_inst|wmgmt_waitrequest[8]~3_combout ;

assign reconfig_mif_address[0] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[0]~q ;

assign reconfig_mif_address[1] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[1]~q ;

assign reconfig_mif_address[2] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[2]~q ;

assign reconfig_mif_address[3] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[3]~q ;

assign reconfig_mif_address[4] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[4]~q ;

assign reconfig_mif_address[5] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[5]~q ;

assign reconfig_mif_address[6] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[6]~q ;

assign reconfig_mif_address[7] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[7]~q ;

assign reconfig_mif_address[8] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[8]~q ;

assign reconfig_mif_address[9] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[9]~q ;

assign reconfig_mif_address[10] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[10]~q ;

assign reconfig_mif_address[11] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[11]~q ;

assign reconfig_mif_address[12] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[12]~q ;

assign reconfig_mif_address[13] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[13]~q ;

assign reconfig_mif_address[14] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[14]~q ;

assign reconfig_mif_address[15] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[15]~q ;

assign reconfig_mif_address[16] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[16]~q ;

assign reconfig_mif_address[17] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[17]~q ;

assign reconfig_mif_address[18] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[18]~q ;

assign reconfig_mif_address[19] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[19]~q ;

assign reconfig_mif_address[20] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[20]~q ;

assign reconfig_mif_address[21] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[21]~q ;

assign reconfig_mif_address[22] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[22]~q ;

assign reconfig_mif_address[23] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[23]~q ;

assign reconfig_mif_address[24] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[24]~q ;

assign reconfig_mif_address[25] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[25]~q ;

assign reconfig_mif_address[26] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[26]~q ;

assign reconfig_mif_address[27] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[27]~q ;

assign reconfig_mif_address[28] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[28]~q ;

assign reconfig_mif_address[29] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[29]~q ;

assign reconfig_mif_address[30] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[30]~q ;

assign reconfig_mif_address[31] = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_address[31]~q ;

assign reconfig_mif_read = \reconfigure_ip_inst|mif.sc_mif|mif_strm_av|inst_mif_avmm|stream_read~q ;

assign reconfig_to_xcvr[0] = \mgmt_clk_clk~input_o ;

assign reconfig_to_xcvr[1] = ~ \reconfigure_ip_inst|inst_reconfig_reset_sync|resync_chains[0].sync_r[1]~q ;

assign reconfig_to_xcvr[2] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[0]~0_combout ;

assign reconfig_to_xcvr[3] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[1]~1_combout ;

assign reconfig_to_xcvr[4] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[2]~2_combout ;

assign reconfig_to_xcvr[5] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[3]~3_combout ;

assign reconfig_to_xcvr[6] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[4]~4_combout ;

assign reconfig_to_xcvr[7] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[5]~5_combout ;

assign reconfig_to_xcvr[8] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[6]~6_combout ;

assign reconfig_to_xcvr[9] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[7]~7_combout ;

assign reconfig_to_xcvr[10] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[8]~8_combout ;

assign reconfig_to_xcvr[11] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[9]~9_combout ;

assign reconfig_to_xcvr[12] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[10]~10_combout ;

assign reconfig_to_xcvr[13] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[11]~11_combout ;

assign reconfig_to_xcvr[14] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[12]~12_combout ;

assign reconfig_to_xcvr[15] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[13]~13_combout ;

assign reconfig_to_xcvr[16] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[14]~14_combout ;

assign reconfig_to_xcvr[17] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[15]~15_combout ;

assign reconfig_to_xcvr[18] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_write[0]~combout ;

assign reconfig_to_xcvr[19] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_read[0]~0_combout ;

assign reconfig_to_xcvr[20] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[0]~combout ;

assign reconfig_to_xcvr[21] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[1]~combout ;

assign reconfig_to_xcvr[22] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[2]~combout ;

assign reconfig_to_xcvr[23] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[3]~combout ;

assign reconfig_to_xcvr[24] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[4]~combout ;

assign reconfig_to_xcvr[25] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[5]~combout ;

assign reconfig_to_xcvr[26] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[6]~combout ;

assign reconfig_to_xcvr[27] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[7]~combout ;

assign reconfig_to_xcvr[28] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[8]~combout ;

assign reconfig_to_xcvr[29] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[9]~combout ;

assign reconfig_to_xcvr[30] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[10]~combout ;

assign reconfig_to_xcvr[31] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[11]~0_combout ;

assign reconfig_to_xcvr[32] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[0]~combout ;

assign reconfig_to_xcvr[33] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[1]~combout ;

assign reconfig_to_xcvr[34] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[2]~combout ;

assign reconfig_to_xcvr[35] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[3]~combout ;

assign reconfig_to_xcvr[36] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[0]~combout ;

assign reconfig_to_xcvr[37] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[1]~combout ;

assign reconfig_to_xcvr[38] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[2]~combout ;

assign reconfig_to_xcvr[39] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[3]~combout ;

assign reconfig_to_xcvr[40] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[0]~combout ;

assign reconfig_to_xcvr[41] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[1]~combout ;

assign reconfig_to_xcvr[42] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[2]~combout ;

assign reconfig_to_xcvr[43] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[3]~combout ;

assign reconfig_to_xcvr[44] = ~ \reconfigure_ip_inst|basic|a5|pif_interface_sel~q ;

assign reconfig_to_xcvr[45] = ~ \reconfigure_ip_inst|basic|a5|pif_ser_shift_load~q ;

assign reconfig_to_xcvr[46] = ~ \reconfigure_ip_inst|offset.sc_offset|offset_cancellation_av|offset_cancellation_done~1_combout ;

assign reconfig_to_xcvr[47] = ~ \reconfigure_ip_inst|cal_seq|tx_cal_busy~q ;

assign reconfig_to_xcvr[48] = ~ \reconfigure_ip_inst|cal_seq|rx_cal_busy~q ;

assign reconfig_to_xcvr[49] = gnd;

assign reconfig_to_xcvr[50] = gnd;

assign reconfig_to_xcvr[51] = gnd;

assign reconfig_to_xcvr[52] = gnd;

assign reconfig_to_xcvr[53] = gnd;

assign reconfig_to_xcvr[54] = gnd;

assign reconfig_to_xcvr[55] = gnd;

assign reconfig_to_xcvr[56] = gnd;

assign reconfig_to_xcvr[57] = gnd;

assign reconfig_to_xcvr[58] = gnd;

assign reconfig_to_xcvr[59] = gnd;

assign reconfig_to_xcvr[60] = gnd;

assign reconfig_to_xcvr[61] = gnd;

assign reconfig_to_xcvr[62] = gnd;

assign reconfig_to_xcvr[63] = gnd;

assign reconfig_to_xcvr[64] = gnd;

assign reconfig_to_xcvr[65] = gnd;

assign reconfig_to_xcvr[66] = gnd;

assign reconfig_to_xcvr[67] = gnd;

assign reconfig_to_xcvr[68] = gnd;

assign reconfig_to_xcvr[69] = gnd;

assign reconfig_to_xcvr[70] = \mgmt_clk_clk~input_o ;

assign reconfig_to_xcvr[71] = ~ \reconfigure_ip_inst|inst_reconfig_reset_sync|resync_chains[0].sync_r[1]~q ;

assign reconfig_to_xcvr[72] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[16]~16_combout ;

assign reconfig_to_xcvr[73] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[17]~17_combout ;

assign reconfig_to_xcvr[74] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[18]~18_combout ;

assign reconfig_to_xcvr[75] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[19]~19_combout ;

assign reconfig_to_xcvr[76] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[20]~20_combout ;

assign reconfig_to_xcvr[77] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[21]~21_combout ;

assign reconfig_to_xcvr[78] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[22]~22_combout ;

assign reconfig_to_xcvr[79] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[23]~23_combout ;

assign reconfig_to_xcvr[80] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[24]~24_combout ;

assign reconfig_to_xcvr[81] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[25]~25_combout ;

assign reconfig_to_xcvr[82] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[26]~26_combout ;

assign reconfig_to_xcvr[83] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[27]~27_combout ;

assign reconfig_to_xcvr[84] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[28]~28_combout ;

assign reconfig_to_xcvr[85] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[29]~29_combout ;

assign reconfig_to_xcvr[86] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[30]~30_combout ;

assign reconfig_to_xcvr[87] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_writedata[31]~31_combout ;

assign reconfig_to_xcvr[88] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_write[1]~combout ;

assign reconfig_to_xcvr[89] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_read[1]~1_combout ;

assign reconfig_to_xcvr[90] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[12]~combout ;

assign reconfig_to_xcvr[91] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[13]~combout ;

assign reconfig_to_xcvr[92] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[14]~combout ;

assign reconfig_to_xcvr[93] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[15]~combout ;

assign reconfig_to_xcvr[94] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[16]~combout ;

assign reconfig_to_xcvr[95] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[17]~combout ;

assign reconfig_to_xcvr[96] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[18]~combout ;

assign reconfig_to_xcvr[97] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[19]~combout ;

assign reconfig_to_xcvr[98] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[20]~combout ;

assign reconfig_to_xcvr[99] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[21]~combout ;

assign reconfig_to_xcvr[100] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[22]~combout ;

assign reconfig_to_xcvr[101] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|native_reconfig_address[23]~1_combout ;

assign reconfig_to_xcvr[102] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[12]~combout ;

assign reconfig_to_xcvr[103] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[13]~combout ;

assign reconfig_to_xcvr[104] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[14]~combout ;

assign reconfig_to_xcvr[105] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[15]~combout ;

assign reconfig_to_xcvr[106] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[12]~combout ;

assign reconfig_to_xcvr[107] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[13]~combout ;

assign reconfig_to_xcvr[108] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[14]~combout ;

assign reconfig_to_xcvr[109] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[15]~combout ;

assign reconfig_to_xcvr[110] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[12]~combout ;

assign reconfig_to_xcvr[111] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[13]~combout ;

assign reconfig_to_xcvr[112] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[14]~combout ;

assign reconfig_to_xcvr[113] = \reconfigure_ip_inst|basic|a5|lif[0].logical_if|pif_testbus_sel[15]~combout ;

assign reconfig_to_xcvr[114] = ~ \reconfigure_ip_inst|basic|a5|pif_interface_sel~q ;

assign reconfig_to_xcvr[115] = ~ \reconfigure_ip_inst|basic|a5|pif_ser_shift_load~q ;

assign reconfig_to_xcvr[116] = ~ \reconfigure_ip_inst|offset.sc_offset|offset_cancellation_av|offset_cancellation_done~1_combout ;

assign reconfig_to_xcvr[117] = ~ \reconfigure_ip_inst|cal_seq|tx_cal_busy~q ;

assign reconfig_to_xcvr[118] = ~ \reconfigure_ip_inst|cal_seq|rx_cal_busy~q ;

assign reconfig_to_xcvr[119] = gnd;

assign reconfig_to_xcvr[120] = gnd;

assign reconfig_to_xcvr[121] = gnd;

assign reconfig_to_xcvr[122] = gnd;

assign reconfig_to_xcvr[123] = gnd;

assign reconfig_to_xcvr[124] = gnd;

assign reconfig_to_xcvr[125] = gnd;

assign reconfig_to_xcvr[126] = gnd;

assign reconfig_to_xcvr[127] = gnd;

assign reconfig_to_xcvr[128] = gnd;

assign reconfig_to_xcvr[129] = gnd;

assign reconfig_to_xcvr[130] = gnd;

assign reconfig_to_xcvr[131] = gnd;

assign reconfig_to_xcvr[132] = gnd;

assign reconfig_to_xcvr[133] = gnd;

assign reconfig_to_xcvr[134] = gnd;

assign reconfig_to_xcvr[135] = gnd;

assign reconfig_to_xcvr[136] = gnd;

assign reconfig_to_xcvr[137] = gnd;

assign reconfig_to_xcvr[138] = gnd;

assign reconfig_to_xcvr[139] = gnd;

assign \mgmt_clk_clk~input_o  = mgmt_clk_clk;

assign \reconfig_from_xcvr[20]~input_o  = reconfig_from_xcvr[20];

assign \reconfig_from_xcvr[21]~input_o  = reconfig_from_xcvr[21];

assign \reconfig_from_xcvr[22]~input_o  = reconfig_from_xcvr[22];

assign \reconfig_from_xcvr[23]~input_o  = reconfig_from_xcvr[23];

assign \reconfig_from_xcvr[28]~input_o  = reconfig_from_xcvr[28];

assign \reconfig_from_xcvr[29]~input_o  = reconfig_from_xcvr[29];

assign \reconfig_from_xcvr[30]~input_o  = reconfig_from_xcvr[30];

assign \reconfig_from_xcvr[31]~input_o  = reconfig_from_xcvr[31];

assign \reconfig_from_xcvr[36]~input_o  = reconfig_from_xcvr[36];

assign \reconfig_from_xcvr[37]~input_o  = reconfig_from_xcvr[37];

assign \reconfig_from_xcvr[38]~input_o  = reconfig_from_xcvr[38];

assign \reconfig_from_xcvr[39]~input_o  = reconfig_from_xcvr[39];

assign \reconfig_from_xcvr[40]~input_o  = reconfig_from_xcvr[40];

assign \reconfig_from_xcvr[41]~input_o  = reconfig_from_xcvr[41];

assign \reconfig_from_xcvr[42]~input_o  = reconfig_from_xcvr[42];

assign \reconfig_from_xcvr[43]~input_o  = reconfig_from_xcvr[43];

assign \reconfig_from_xcvr[44]~input_o  = reconfig_from_xcvr[44];

assign \reconfig_from_xcvr[45]~input_o  = reconfig_from_xcvr[45];

assign \reconfig_from_xcvr[66]~input_o  = reconfig_from_xcvr[66];

assign \reconfig_from_xcvr[67]~input_o  = reconfig_from_xcvr[67];

assign \reconfig_from_xcvr[68]~input_o  = reconfig_from_xcvr[68];

assign \reconfig_from_xcvr[69]~input_o  = reconfig_from_xcvr[69];

assign \reconfig_from_xcvr[74]~input_o  = reconfig_from_xcvr[74];

assign \reconfig_from_xcvr[75]~input_o  = reconfig_from_xcvr[75];

assign \reconfig_from_xcvr[76]~input_o  = reconfig_from_xcvr[76];

assign \reconfig_from_xcvr[77]~input_o  = reconfig_from_xcvr[77];

assign \reconfig_from_xcvr[82]~input_o  = reconfig_from_xcvr[82];

assign \reconfig_from_xcvr[83]~input_o  = reconfig_from_xcvr[83];

assign \reconfig_from_xcvr[84]~input_o  = reconfig_from_xcvr[84];

assign \reconfig_from_xcvr[85]~input_o  = reconfig_from_xcvr[85];

assign \reconfig_from_xcvr[86]~input_o  = reconfig_from_xcvr[86];

assign \reconfig_from_xcvr[87]~input_o  = reconfig_from_xcvr[87];

assign \reconfig_from_xcvr[88]~input_o  = reconfig_from_xcvr[88];

assign \reconfig_from_xcvr[89]~input_o  = reconfig_from_xcvr[89];

assign \reconfig_from_xcvr[90]~input_o  = reconfig_from_xcvr[90];

assign \reconfig_from_xcvr[91]~input_o  = reconfig_from_xcvr[91];

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig (
	stream_address_0,
	stream_address_1,
	stream_address_2,
	stream_address_3,
	stream_address_4,
	stream_address_5,
	stream_address_6,
	stream_address_7,
	stream_address_8,
	stream_address_9,
	stream_address_10,
	stream_address_11,
	stream_address_12,
	stream_address_13,
	stream_address_14,
	stream_address_15,
	stream_address_16,
	stream_address_17,
	stream_address_18,
	stream_address_19,
	stream_address_20,
	stream_address_21,
	stream_address_22,
	stream_address_23,
	stream_address_24,
	stream_address_25,
	stream_address_26,
	stream_address_27,
	stream_address_28,
	stream_address_29,
	stream_address_30,
	stream_address_31,
	rtl,
	reconfig_busy,
	wmgmt_readdata_0_8,
	wmgmt_readdata_1_8,
	wmgmt_readdata_2_8,
	wmgmt_readdata_3_8,
	wmgmt_readdata_4_8,
	wmgmt_readdata_5_8,
	wmgmt_readdata_6_8,
	wmgmt_readdata_7_8,
	reconfig_mgmt_readdata_8,
	wmgmt_readdata_9_8,
	wmgmt_readdata_10_8,
	wmgmt_readdata_11_8,
	wmgmt_readdata_12_8,
	wmgmt_readdata_13_8,
	wmgmt_readdata_14_8,
	wmgmt_readdata_15_8,
	wmgmt_readdata_16_8,
	wmgmt_readdata_17_8,
	wmgmt_readdata_18_8,
	wmgmt_readdata_19_8,
	wmgmt_readdata_20_8,
	wmgmt_readdata_21_8,
	wmgmt_readdata_22_8,
	wmgmt_readdata_23_8,
	wmgmt_readdata_24_8,
	wmgmt_readdata_25_8,
	wmgmt_readdata_26_8,
	wmgmt_readdata_27_8,
	wmgmt_readdata_28_8,
	wmgmt_readdata_29_8,
	wmgmt_readdata_30_8,
	wmgmt_readdata_31_8,
	wmgmt_waitrequest_8,
	stream_read,
	resync_chains0sync_r_1,
	native_reconfig_writedata_0,
	native_reconfig_writedata_1,
	native_reconfig_writedata_2,
	native_reconfig_writedata_3,
	native_reconfig_writedata_4,
	native_reconfig_writedata_5,
	native_reconfig_writedata_6,
	native_reconfig_writedata_7,
	native_reconfig_writedata_8,
	native_reconfig_writedata_9,
	native_reconfig_writedata_10,
	native_reconfig_writedata_11,
	native_reconfig_writedata_12,
	native_reconfig_writedata_13,
	native_reconfig_writedata_14,
	native_reconfig_writedata_15,
	native_reconfig_write_0,
	native_reconfig_read_0,
	native_reconfig_address_0,
	native_reconfig_address_1,
	native_reconfig_address_2,
	native_reconfig_address_3,
	native_reconfig_address_4,
	native_reconfig_address_5,
	native_reconfig_address_6,
	native_reconfig_address_7,
	native_reconfig_address_8,
	native_reconfig_address_9,
	native_reconfig_address_10,
	native_reconfig_address_11,
	pif_testbus_sel_0,
	pif_testbus_sel_1,
	pif_testbus_sel_2,
	pif_testbus_sel_3,
	pif_interface_sel,
	pif_ser_shift_load,
	offset_cancellation_done,
	tx_cal_busy,
	rx_cal_busy,
	native_reconfig_writedata_16,
	native_reconfig_writedata_17,
	native_reconfig_writedata_18,
	native_reconfig_writedata_19,
	native_reconfig_writedata_20,
	native_reconfig_writedata_21,
	native_reconfig_writedata_22,
	native_reconfig_writedata_23,
	native_reconfig_writedata_24,
	native_reconfig_writedata_25,
	native_reconfig_writedata_26,
	native_reconfig_writedata_27,
	native_reconfig_writedata_28,
	native_reconfig_writedata_29,
	native_reconfig_writedata_30,
	native_reconfig_writedata_31,
	native_reconfig_write_1,
	native_reconfig_read_1,
	native_reconfig_address_12,
	native_reconfig_address_13,
	native_reconfig_address_14,
	native_reconfig_address_15,
	native_reconfig_address_16,
	native_reconfig_address_17,
	native_reconfig_address_18,
	native_reconfig_address_19,
	native_reconfig_address_20,
	native_reconfig_address_21,
	native_reconfig_address_22,
	native_reconfig_address_23,
	pif_testbus_sel_12,
	pif_testbus_sel_13,
	pif_testbus_sel_14,
	pif_testbus_sel_15,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_0,
	Decoder3,
	readdata_for_user_2,
	readdata_for_user_0,
	readdata_for_user_3,
	readdata_for_user_1,
	Decoder31,
	Selector2,
	Selector21,
	Decoder32,
	lpbk_lock,
	analog_offset_0,
	readdata_for_user_10,
	readdata_for_user_8,
	readdata_for_user_11,
	readdata_for_user_9,
	rtl1,
	readdata_for_user_6,
	readdata_for_user_4,
	readdata_for_user_7,
	readdata_for_user_5,
	readdata_for_user_14,
	readdata_for_user_12,
	readdata_for_user_15,
	readdata_for_user_13,
	rtl2,
	rtl3,
	rtl4,
	rtl5,
	rtl6,
	readdata_for_user_16,
	rtl7,
	rtl8,
	WideOr4,
	WideOr41,
	analog_length,
	analog_length1,
	analog_length2,
	rtl9,
	readdata_for_user_17,
	rtl10,
	rtl11,
	rtl12,
	readdata_for_user_18,
	rtl13,
	rtl14,
	uif_writedata_4,
	readdata_for_user_19,
	rtl15,
	rtl16,
	LessThan4,
	readdata_for_user_20,
	rtl17,
	rtl18,
	readdata_for_user_21,
	rtl19,
	rtl20,
	readdata_for_user_22,
	rtl21,
	rtl22,
	readdata_for_user_23,
	rtl23,
	readdata_for_user_24,
	rtl24,
	readdata_for_user_25,
	rtl25,
	readdata_for_user_26,
	rtl26,
	readdata_for_user_27,
	rtl27,
	readdata_for_user_28,
	rtl28,
	readdata_for_user_29,
	rtl29,
	readdata_for_user_30,
	rtl30,
	readdata_for_user_31,
	rtl31,
	rtl32,
	rtl33,
	Selector5,
	result_data_0,
	rtl34,
	rtl35,
	rtl36,
	rtl37,
	rtl38,
	rtl39,
	rtl40,
	rtl41,
	rtl42,
	rtl43,
	GND_port,
	reconfig_mgmt_address_3,
	reconfig_mgmt_address_4,
	reconfig_mgmt_address_5,
	reconfig_mgmt_address_6,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mif_waitrequest,
	reconfig_mgmt_writedata_16,
	reconfig_from_xcvr_0,
	reconfig_from_xcvr_46,
	reconfig_mgmt_writedata_17,
	reconfig_from_xcvr_1,
	reconfig_from_xcvr_47,
	reconfig_mgmt_writedata_18,
	reconfig_from_xcvr_2,
	reconfig_from_xcvr_48,
	reconfig_mgmt_writedata_19,
	reconfig_from_xcvr_3,
	reconfig_from_xcvr_49,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_from_xcvr_4,
	reconfig_from_xcvr_50,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_from_xcvr_5,
	reconfig_from_xcvr_51,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_from_xcvr_6,
	reconfig_from_xcvr_52,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_from_xcvr_7,
	reconfig_from_xcvr_53,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_from_xcvr_8,
	reconfig_from_xcvr_54,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_from_xcvr_9,
	reconfig_from_xcvr_55,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_from_xcvr_10,
	reconfig_from_xcvr_56,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_from_xcvr_11,
	reconfig_from_xcvr_57,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_from_xcvr_12,
	reconfig_from_xcvr_58,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_from_xcvr_13,
	reconfig_from_xcvr_59,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_from_xcvr_14,
	reconfig_from_xcvr_60,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15,
	reconfig_from_xcvr_15,
	reconfig_from_xcvr_61,
	reconfig_mif_readdata_15,
	reconfig_mif_readdata_14,
	reconfig_mif_readdata_13,
	reconfig_mif_readdata_12,
	reconfig_mif_readdata_11,
	reconfig_mif_readdata_1,
	reconfig_mif_readdata_0,
	reconfig_mif_readdata_4,
	reconfig_mif_readdata_3,
	reconfig_mif_readdata_2,
	mgmt_rst_reset,
	reconfig_mif_readdata_7,
	reconfig_mif_readdata_5,
	reconfig_mif_readdata_6,
	reconfig_mif_readdata_8,
	reconfig_mif_readdata_9,
	reconfig_mif_readdata_10,
	reconfig_from_xcvr_24,
	reconfig_from_xcvr_70,
	reconfig_from_xcvr_16,
	reconfig_from_xcvr_62,
	reconfig_from_xcvr_32,
	reconfig_from_xcvr_78,
	reconfig_from_xcvr_25,
	reconfig_from_xcvr_71,
	reconfig_from_xcvr_17,
	reconfig_from_xcvr_63,
	reconfig_from_xcvr_33,
	reconfig_from_xcvr_79,
	reconfig_from_xcvr_26,
	reconfig_from_xcvr_72,
	reconfig_from_xcvr_18,
	reconfig_from_xcvr_64,
	reconfig_from_xcvr_34,
	reconfig_from_xcvr_80,
	reconfig_from_xcvr_27,
	reconfig_from_xcvr_73,
	reconfig_from_xcvr_19,
	reconfig_from_xcvr_65,
	reconfig_from_xcvr_35,
	reconfig_from_xcvr_81)/* synthesis synthesis_greybox=0 */;
output 	stream_address_0;
output 	stream_address_1;
output 	stream_address_2;
output 	stream_address_3;
output 	stream_address_4;
output 	stream_address_5;
output 	stream_address_6;
output 	stream_address_7;
output 	stream_address_8;
output 	stream_address_9;
output 	stream_address_10;
output 	stream_address_11;
output 	stream_address_12;
output 	stream_address_13;
output 	stream_address_14;
output 	stream_address_15;
output 	stream_address_16;
output 	stream_address_17;
output 	stream_address_18;
output 	stream_address_19;
output 	stream_address_20;
output 	stream_address_21;
output 	stream_address_22;
output 	stream_address_23;
output 	stream_address_24;
output 	stream_address_25;
output 	stream_address_26;
output 	stream_address_27;
output 	stream_address_28;
output 	stream_address_29;
output 	stream_address_30;
output 	stream_address_31;
input 	rtl;
output 	reconfig_busy;
output 	wmgmt_readdata_0_8;
output 	wmgmt_readdata_1_8;
output 	wmgmt_readdata_2_8;
output 	wmgmt_readdata_3_8;
output 	wmgmt_readdata_4_8;
output 	wmgmt_readdata_5_8;
output 	wmgmt_readdata_6_8;
output 	wmgmt_readdata_7_8;
output 	reconfig_mgmt_readdata_8;
output 	wmgmt_readdata_9_8;
output 	wmgmt_readdata_10_8;
output 	wmgmt_readdata_11_8;
output 	wmgmt_readdata_12_8;
output 	wmgmt_readdata_13_8;
output 	wmgmt_readdata_14_8;
output 	wmgmt_readdata_15_8;
output 	wmgmt_readdata_16_8;
output 	wmgmt_readdata_17_8;
output 	wmgmt_readdata_18_8;
output 	wmgmt_readdata_19_8;
output 	wmgmt_readdata_20_8;
output 	wmgmt_readdata_21_8;
output 	wmgmt_readdata_22_8;
output 	wmgmt_readdata_23_8;
output 	wmgmt_readdata_24_8;
output 	wmgmt_readdata_25_8;
output 	wmgmt_readdata_26_8;
output 	wmgmt_readdata_27_8;
output 	wmgmt_readdata_28_8;
output 	wmgmt_readdata_29_8;
output 	wmgmt_readdata_30_8;
output 	wmgmt_readdata_31_8;
output 	wmgmt_waitrequest_8;
output 	stream_read;
output 	resync_chains0sync_r_1;
output 	native_reconfig_writedata_0;
output 	native_reconfig_writedata_1;
output 	native_reconfig_writedata_2;
output 	native_reconfig_writedata_3;
output 	native_reconfig_writedata_4;
output 	native_reconfig_writedata_5;
output 	native_reconfig_writedata_6;
output 	native_reconfig_writedata_7;
output 	native_reconfig_writedata_8;
output 	native_reconfig_writedata_9;
output 	native_reconfig_writedata_10;
output 	native_reconfig_writedata_11;
output 	native_reconfig_writedata_12;
output 	native_reconfig_writedata_13;
output 	native_reconfig_writedata_14;
output 	native_reconfig_writedata_15;
output 	native_reconfig_write_0;
output 	native_reconfig_read_0;
output 	native_reconfig_address_0;
output 	native_reconfig_address_1;
output 	native_reconfig_address_2;
output 	native_reconfig_address_3;
output 	native_reconfig_address_4;
output 	native_reconfig_address_5;
output 	native_reconfig_address_6;
output 	native_reconfig_address_7;
output 	native_reconfig_address_8;
output 	native_reconfig_address_9;
output 	native_reconfig_address_10;
output 	native_reconfig_address_11;
output 	pif_testbus_sel_0;
output 	pif_testbus_sel_1;
output 	pif_testbus_sel_2;
output 	pif_testbus_sel_3;
output 	pif_interface_sel;
output 	pif_ser_shift_load;
output 	offset_cancellation_done;
output 	tx_cal_busy;
output 	rx_cal_busy;
output 	native_reconfig_writedata_16;
output 	native_reconfig_writedata_17;
output 	native_reconfig_writedata_18;
output 	native_reconfig_writedata_19;
output 	native_reconfig_writedata_20;
output 	native_reconfig_writedata_21;
output 	native_reconfig_writedata_22;
output 	native_reconfig_writedata_23;
output 	native_reconfig_writedata_24;
output 	native_reconfig_writedata_25;
output 	native_reconfig_writedata_26;
output 	native_reconfig_writedata_27;
output 	native_reconfig_writedata_28;
output 	native_reconfig_writedata_29;
output 	native_reconfig_writedata_30;
output 	native_reconfig_writedata_31;
output 	native_reconfig_write_1;
output 	native_reconfig_read_1;
output 	native_reconfig_address_12;
output 	native_reconfig_address_13;
output 	native_reconfig_address_14;
output 	native_reconfig_address_15;
output 	native_reconfig_address_16;
output 	native_reconfig_address_17;
output 	native_reconfig_address_18;
output 	native_reconfig_address_19;
output 	native_reconfig_address_20;
output 	native_reconfig_address_21;
output 	native_reconfig_address_22;
output 	native_reconfig_address_23;
output 	pif_testbus_sel_12;
output 	pif_testbus_sel_13;
output 	pif_testbus_sel_14;
output 	pif_testbus_sel_15;
output 	uif_addr_offset_5;
output 	uif_addr_offset_4;
output 	uif_addr_offset_0;
output 	Decoder3;
output 	readdata_for_user_2;
output 	readdata_for_user_0;
output 	readdata_for_user_3;
output 	readdata_for_user_1;
output 	Decoder31;
output 	Selector2;
output 	Selector21;
output 	Decoder32;
output 	lpbk_lock;
output 	analog_offset_0;
output 	readdata_for_user_10;
output 	readdata_for_user_8;
output 	readdata_for_user_11;
output 	readdata_for_user_9;
input 	rtl1;
output 	readdata_for_user_6;
output 	readdata_for_user_4;
output 	readdata_for_user_7;
output 	readdata_for_user_5;
output 	readdata_for_user_14;
output 	readdata_for_user_12;
output 	readdata_for_user_15;
output 	readdata_for_user_13;
input 	rtl2;
input 	rtl3;
input 	rtl4;
input 	rtl5;
input 	rtl6;
output 	readdata_for_user_16;
input 	rtl7;
input 	rtl8;
output 	WideOr4;
output 	WideOr41;
output 	analog_length;
output 	analog_length1;
output 	analog_length2;
input 	rtl9;
output 	readdata_for_user_17;
input 	rtl10;
input 	rtl11;
input 	rtl12;
output 	readdata_for_user_18;
input 	rtl13;
input 	rtl14;
output 	uif_writedata_4;
output 	readdata_for_user_19;
input 	rtl15;
input 	rtl16;
output 	LessThan4;
output 	readdata_for_user_20;
input 	rtl17;
input 	rtl18;
output 	readdata_for_user_21;
input 	rtl19;
input 	rtl20;
output 	readdata_for_user_22;
input 	rtl21;
input 	rtl22;
output 	readdata_for_user_23;
input 	rtl23;
output 	readdata_for_user_24;
input 	rtl24;
output 	readdata_for_user_25;
input 	rtl25;
output 	readdata_for_user_26;
input 	rtl26;
output 	readdata_for_user_27;
input 	rtl27;
output 	readdata_for_user_28;
input 	rtl28;
output 	readdata_for_user_29;
input 	rtl29;
output 	readdata_for_user_30;
input 	rtl30;
output 	readdata_for_user_31;
input 	rtl31;
input 	rtl32;
input 	rtl33;
output 	Selector5;
output 	result_data_0;
input 	rtl34;
input 	rtl35;
input 	rtl36;
input 	rtl37;
input 	rtl38;
input 	rtl39;
input 	rtl40;
input 	rtl41;
input 	rtl42;
input 	rtl43;
input 	GND_port;
input 	reconfig_mgmt_address_3;
input 	reconfig_mgmt_address_4;
input 	reconfig_mgmt_address_5;
input 	reconfig_mgmt_address_6;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mif_waitrequest;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_from_xcvr_0;
input 	reconfig_from_xcvr_46;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_from_xcvr_1;
input 	reconfig_from_xcvr_47;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_from_xcvr_2;
input 	reconfig_from_xcvr_48;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_from_xcvr_3;
input 	reconfig_from_xcvr_49;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_from_xcvr_4;
input 	reconfig_from_xcvr_50;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_from_xcvr_5;
input 	reconfig_from_xcvr_51;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_from_xcvr_6;
input 	reconfig_from_xcvr_52;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_from_xcvr_7;
input 	reconfig_from_xcvr_53;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_from_xcvr_8;
input 	reconfig_from_xcvr_54;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_from_xcvr_9;
input 	reconfig_from_xcvr_55;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_from_xcvr_10;
input 	reconfig_from_xcvr_56;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_from_xcvr_11;
input 	reconfig_from_xcvr_57;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_from_xcvr_12;
input 	reconfig_from_xcvr_58;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_from_xcvr_13;
input 	reconfig_from_xcvr_59;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_from_xcvr_14;
input 	reconfig_from_xcvr_60;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;
input 	reconfig_from_xcvr_15;
input 	reconfig_from_xcvr_61;
input 	reconfig_mif_readdata_15;
input 	reconfig_mif_readdata_14;
input 	reconfig_mif_readdata_13;
input 	reconfig_mif_readdata_12;
input 	reconfig_mif_readdata_11;
input 	reconfig_mif_readdata_1;
input 	reconfig_mif_readdata_0;
input 	reconfig_mif_readdata_4;
input 	reconfig_mif_readdata_3;
input 	reconfig_mif_readdata_2;
input 	mgmt_rst_reset;
input 	reconfig_mif_readdata_7;
input 	reconfig_mif_readdata_5;
input 	reconfig_mif_readdata_6;
input 	reconfig_mif_readdata_8;
input 	reconfig_mif_readdata_9;
input 	reconfig_mif_readdata_10;
input 	reconfig_from_xcvr_24;
input 	reconfig_from_xcvr_70;
input 	reconfig_from_xcvr_16;
input 	reconfig_from_xcvr_62;
input 	reconfig_from_xcvr_32;
input 	reconfig_from_xcvr_78;
input 	reconfig_from_xcvr_25;
input 	reconfig_from_xcvr_71;
input 	reconfig_from_xcvr_17;
input 	reconfig_from_xcvr_63;
input 	reconfig_from_xcvr_33;
input 	reconfig_from_xcvr_79;
input 	reconfig_from_xcvr_26;
input 	reconfig_from_xcvr_72;
input 	reconfig_from_xcvr_18;
input 	reconfig_from_xcvr_64;
input 	reconfig_from_xcvr_34;
input 	reconfig_from_xcvr_80;
input 	reconfig_from_xcvr_27;
input 	reconfig_from_xcvr_73;
input 	reconfig_from_xcvr_19;
input 	reconfig_from_xcvr_65;
input 	reconfig_from_xcvr_35;
input 	reconfig_from_xcvr_81;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[6]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[7]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[10]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[10]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[11]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[11]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[12]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[12]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[12]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[12]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[13]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[13]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[13]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[13]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[14]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[14]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[14]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[14]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[15]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[15]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[15]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[15]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[16]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[16]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[16]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[16]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[17]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[17]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[17]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[17]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[18]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[18]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[18]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[18]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[19]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[19]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[19]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[19]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[20]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[20]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[20]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[21]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[21]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[21]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[22]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[22]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[22]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[23]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[23]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[23]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[24]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[24]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[24]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[25]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[25]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[26]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[26]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[27]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[27]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[28]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[28]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[29]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[29]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[30]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[30]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[31]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[31]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[16]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[17]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[18]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[19]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[20]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[21]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[22]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[23]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[24]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[25]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[26]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[27]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[28]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[29]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[30]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[31]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[0]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[0]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[0]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[0]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[1]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[1]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[1]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[1]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[2]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[2]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[2]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[2]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[3]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[3]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[3]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[3]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[4]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[4]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[4]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[4]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[5]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[5]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[5]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[5]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[6]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[6]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[6]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[7]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[7]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[7]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[8]~q ;
wire \offset.sc_offset|offset_cancellation_av|offset_cancellation_readdata[8]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[8]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[8]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[8]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[9]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[9]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[9]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[9]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[10]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[10]~q ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[11]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[11]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[20]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[21]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[22]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[23]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[24]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[25]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[25]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[26]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[26]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[27]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[27]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[28]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[28]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[29]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[29]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[30]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[30]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[31]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[31]~q ;
wire \direct.sc_direct|reg_arb_req~q ;
wire \arbiter|grant[4]~q ;
wire \direct.sc_direct|mutex_inst|mutex_grant~combout ;
wire \direct.sc_direct|mutex_inst|master_write~0_combout ;
wire \offset.sc_offset|offset_cancellation_av|master_write~q ;
wire \arbiter|grant[0]~q ;
wire \offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_write~q ;
wire \arbiter|grant[1]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ;
wire \wbasic_write[8]~0_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_write~q ;
wire \arbiter|grant[7]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_write~q ;
wire \arbiter|grant[8]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ;
wire \wbasic_write[8]~1_combout ;
wire \wbasic_write[8]~2_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[2]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_address[2]~combout ;
wire \offset.sc_offset|offset_cancellation_av|master_address[2]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[2]~q ;
wire \wbasic_address[8][2]~0_combout ;
wire \wbasic_address[8][2]~combout ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_address[0]~q ;
wire \wbasic_address[8][0]~1_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ;
wire \wbasic_address[8][0]~2_combout ;
wire \wbasic_address[8][0]~3_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[1]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_address[1]~combout ;
wire \offset.sc_offset|offset_cancellation_av|master_address[1]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[1]~q ;
wire \wbasic_address[8][1]~4_combout ;
wire \wbasic_address[8][1]~combout ;
wire \basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~1_combout ;
wire \offset.sc_offset|offset_cancellation_av|master_read~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_read~q ;
wire \wbasic_read[8]~0_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_read~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_read~q ;
wire \wbasic_read[8]~1_combout ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~0_combout ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~1_combout ;
wire \offset.sc_offset|offset_cancellation_av|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ;
wire \offset.sc_offset|offset_cancellation_av|wait_gen|launch_reg~q ;
wire \offset.sc_offset|offset_cancellation_av|wait_gen|wait_reg~q ;
wire \comb~0_combout ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|wait_gen|wait_req~0_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|launch_reg~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|wait_reg~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|launch_reg~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|wait_reg~q ;
wire \mif.sc_mif|mif_strm_av|inst_mif_ctrl|uif_busy~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_ctrl|pll_mif_busy~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|inst_analog_ctrlsm|state.STATE_IDLE~q ;
wire \ifsel_notdone_resync~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[0]~q ;
wire \comb~1_combout ;
wire \comb~2_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[1]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[2]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[3]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[10]~7_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[4]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[5]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[6]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[7]~q ;
wire \comb~3_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[8]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[9]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ;
wire \arbiter|WideNor0~combout ;
wire \offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ;
wire \basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~5_combout ;
wire \direct.sc_direct|mutex_inst|master_read~combout ;
wire \wbasic_read[8]~2_combout ;
wire \basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~6_combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|Equal8~0_combout ;
wire \basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~2_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[1]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[1]~combout ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[1]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[1]~q ;
wire \wbasic_writedata[8][1]~0_combout ;
wire \wbasic_writedata[8][1]~combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[2]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[2]~combout ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[2]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[2]~q ;
wire \wbasic_writedata[8][2]~1_combout ;
wire \wbasic_writedata[8][2]~combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[0]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[0]~combout ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[0]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[0]~q ;
wire \wbasic_writedata[8][0]~2_combout ;
wire \wbasic_writedata[8][0]~combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[3]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[3]~combout ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[3]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[3]~q ;
wire \wbasic_writedata[8][3]~3_combout ;
wire \wbasic_writedata[8][3]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[4]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ;
wire \wbasic_writedata[8][4]~4_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ;
wire \wbasic_writedata[8][4]~5_combout ;
wire \wbasic_writedata[8][4]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[5]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ;
wire \wbasic_writedata[8][5]~6_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ;
wire \wbasic_writedata[8][5]~7_combout ;
wire \wbasic_writedata[8][5]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[6]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ;
wire \wbasic_writedata[8][6]~8_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ;
wire \wbasic_writedata[8][6]~9_combout ;
wire \wbasic_writedata[8][6]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[7]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ;
wire \wbasic_writedata[8][7]~10_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ;
wire \wbasic_writedata[8][7]~11_combout ;
wire \wbasic_writedata[8][7]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[8]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ;
wire \wbasic_writedata[8][8]~12_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ;
wire \wbasic_writedata[8][8]~13_combout ;
wire \wbasic_writedata[8][8]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[9]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ;
wire \wbasic_writedata[8][9]~14_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ;
wire \wbasic_writedata[8][9]~15_combout ;
wire \wbasic_writedata[8][9]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[10]~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ;
wire \wbasic_writedata[8][10]~16_combout ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ;
wire \wbasic_writedata[8][10]~17_combout ;
wire \wbasic_writedata[8][10]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[11]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ;
wire \wbasic_writedata[8][11]~18_combout ;
wire \wbasic_writedata[8][11]~19_combout ;
wire \wbasic_writedata[8][11]~combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[12]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[13]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[14]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ;
wire \pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ;
wire \offset.sc_offset|offset_cancellation_av|master_write_data[15]~q ;
wire \mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ;
wire \basic|a5|LessThan0~0_combout ;
wire \mif.sc_mif|mif_strm_av|inst_mif_avmm|pll_go~q ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_mode[0]~0_combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux0~0_combout ;
wire \pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux3~0_combout ;
wire \wbasic_write[8]~combout ;
wire \reg_grant_last[4]~q ;
wire \reg_grant_last[7]~q ;
wire \reg_grant_last[8]~q ;
wire \lif_is_active~0_combout ;
wire \reg_grant_last[0]~q ;
wire \reg_grant_last[1]~q ;
wire \lif_is_active~1_combout ;
wire \lif_is_active~combout ;
wire \analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|WideOr0~0_combout ;
wire \mif.sc_mif|mif_strm_av|inst_mif_avmm|pll_type~q ;
wire \mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[7]~q ;
wire \mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[5]~q ;
wire \mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[6]~q ;
wire \basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[0]~combout ;
wire \basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[1]~combout ;
wire \basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[2]~combout ;
wire \basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[3]~combout ;
wire \Equal3~0_combout ;
wire \Equal4~0_combout ;
wire \wmgmt_readdata[8][0]~0_combout ;
wire \wmgmt_readdata[8][1]~1_combout ;
wire \wmgmt_readdata[8][2]~2_combout ;
wire \wmgmt_readdata[8][3]~3_combout ;
wire \wmgmt_readdata[8][4]~4_combout ;
wire \wmgmt_readdata[8][5]~5_combout ;
wire \Equal1~0_combout ;
wire \Equal2~0_combout ;
wire \wmgmt_readdata[8][6]~6_combout ;
wire \wmgmt_readdata[8][7]~7_combout ;
wire \reconfig_mgmt_readdata[8]~0_combout ;
wire \reconfig_mgmt_readdata[8]~1_combout ;
wire \reconfig_mgmt_readdata[8]~2_combout ;
wire \wmgmt_readdata[8][9]~8_combout ;
wire \wmgmt_readdata~9_combout ;
wire \wmgmt_readdata~10_combout ;
wire \wmgmt_readdata~11_combout ;
wire \wmgmt_readdata~12_combout ;
wire \wmgmt_readdata[8][12]~13_combout ;
wire \wmgmt_readdata[8][13]~14_combout ;
wire \wmgmt_readdata[8][14]~15_combout ;
wire \wmgmt_readdata[8][15]~16_combout ;
wire \wmgmt_readdata[8][16]~17_combout ;
wire \wmgmt_readdata[8][17]~18_combout ;
wire \wmgmt_readdata[8][18]~19_combout ;
wire \wmgmt_readdata[8][19]~20_combout ;
wire \wmgmt_readdata[8][20]~21_combout ;
wire \wmgmt_readdata[8][21]~22_combout ;
wire \wmgmt_readdata[8][22]~23_combout ;
wire \wmgmt_readdata[8][23]~24_combout ;
wire \wmgmt_readdata[8][24]~25_combout ;
wire \wmgmt_readdata~26_combout ;
wire \wmgmt_readdata~27_combout ;
wire \wmgmt_readdata~28_combout ;
wire \wmgmt_readdata~29_combout ;
wire \wmgmt_readdata~30_combout ;
wire \wmgmt_readdata~31_combout ;
wire \wmgmt_readdata~32_combout ;
wire \wmgmt_readdata~33_combout ;
wire \wmgmt_readdata~34_combout ;
wire \wmgmt_readdata~35_combout ;
wire \wmgmt_readdata~36_combout ;
wire \wmgmt_readdata~37_combout ;
wire \wmgmt_readdata~38_combout ;
wire \wmgmt_readdata~39_combout ;
wire \Equal0~0_combout ;
wire \wmgmt_waitrequest[0]~combout ;
wire \wmgmt_waitrequest~0_combout ;
wire \wmgmt_waitrequest~1_combout ;
wire \wmgmt_waitrequest[8]~2_combout ;


RECONFIGURE_IP_alt_xcvr_reconfig_offset_cancellation \offset.sc_offset (
	.basic_reconfig_readdata_12(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[12]~q ),
	.basic_reconfig_readdata_13(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[13]~q ),
	.basic_reconfig_readdata_14(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[14]~q ),
	.basic_reconfig_readdata_15(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[15]~q ),
	.basic_reconfig_readdata_0(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[0]~q ),
	.basic_reconfig_readdata_1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[1]~q ),
	.basic_reconfig_readdata_2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[2]~q ),
	.basic_reconfig_readdata_3(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[3]~q ),
	.basic_reconfig_readdata_4(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[4]~q ),
	.basic_reconfig_readdata_5(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[5]~q ),
	.basic_reconfig_readdata_6(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[6]~q ),
	.basic_reconfig_readdata_7(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[7]~q ),
	.reconfig_mgmt_readdata_8(\reconfig_mgmt_readdata[8]~0_combout ),
	.offset_cancellation_readdata_8(\offset.sc_offset|offset_cancellation_av|offset_cancellation_readdata[8]~q ),
	.basic_reconfig_readdata_8(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[8]~q ),
	.basic_reconfig_readdata_9(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_10(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[10]~q ),
	.basic_reconfig_readdata_11(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[11]~q ),
	.master_write(\offset.sc_offset|offset_cancellation_av|master_write~q ),
	.grant_0(\arbiter|grant[0]~q ),
	.req_and_use_mutex(\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.master_address_2(\offset.sc_offset|offset_cancellation_av|master_address[2]~q ),
	.master_address_0(\offset.sc_offset|offset_cancellation_av|master_address[0]~q ),
	.master_address_1(\offset.sc_offset|offset_cancellation_av|master_address[1]~q ),
	.lif_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~1_combout ),
	.master_read(\offset.sc_offset|offset_cancellation_av|master_read~q ),
	.basic_reconfig_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~0_combout ),
	.basic_reconfig_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~1_combout ),
	.Equal0(\Equal0~0_combout ),
	.resync_chains0sync_r_1(\offset.sc_offset|offset_cancellation_av|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ),
	.launch_reg(\offset.sc_offset|offset_cancellation_av|wait_gen|launch_reg~q ),
	.wait_reg(\offset.sc_offset|offset_cancellation_av|wait_gen|wait_reg~q ),
	.offset_cancellation_done(offset_cancellation_done),
	.ifsel_notdone_resync(\ifsel_notdone_resync~q ),
	.comb(\comb~3_combout ),
	.mutex_grant(\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.lif_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~5_combout ),
	.lif_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~6_combout ),
	.Equal8(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|Equal8~0_combout ),
	.basic_reconfig_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~2_combout ),
	.master_write_data_1(\offset.sc_offset|offset_cancellation_av|master_write_data[1]~q ),
	.master_write_data_2(\offset.sc_offset|offset_cancellation_av|master_write_data[2]~q ),
	.master_write_data_0(\offset.sc_offset|offset_cancellation_av|master_write_data[0]~q ),
	.master_write_data_3(\offset.sc_offset|offset_cancellation_av|master_write_data[3]~q ),
	.master_write_data_4(\offset.sc_offset|offset_cancellation_av|master_write_data[4]~q ),
	.master_write_data_5(\offset.sc_offset|offset_cancellation_av|master_write_data[5]~q ),
	.master_write_data_6(\offset.sc_offset|offset_cancellation_av|master_write_data[6]~q ),
	.master_write_data_7(\offset.sc_offset|offset_cancellation_av|master_write_data[7]~q ),
	.master_write_data_8(\offset.sc_offset|offset_cancellation_av|master_write_data[8]~q ),
	.master_write_data_9(\offset.sc_offset|offset_cancellation_av|master_write_data[9]~q ),
	.master_write_data_10(\offset.sc_offset|offset_cancellation_av|master_write_data[10]~q ),
	.master_write_data_11(\offset.sc_offset|offset_cancellation_av|master_write_data[11]~q ),
	.master_write_data_12(\offset.sc_offset|offset_cancellation_av|master_write_data[12]~q ),
	.master_write_data_13(\offset.sc_offset|offset_cancellation_av|master_write_data[13]~q ),
	.master_write_data_14(\offset.sc_offset|offset_cancellation_av|master_write_data[14]~q ),
	.master_write_data_15(\offset.sc_offset|offset_cancellation_av|master_write_data[15]~q ),
	.out_narrow_0(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[0]~combout ),
	.out_narrow_1(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[1]~combout ),
	.out_narrow_2(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[2]~combout ),
	.out_narrow_3(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[3]~combout ),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0));

RECONFIGURE_IP_alt_xcvr_resync_4 inst_reconfig_reset_sync(
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.clk(mgmt_clk_clk),
	.mgmt_rst_reset(mgmt_rst_reset));

RECONFIGURE_IP_alt_xcvr_arbiter arbiter(
	.reg_arb_req(\direct.sc_direct|reg_arb_req~q ),
	.grant_4(\arbiter|grant[4]~q ),
	.mutex_grant(\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.grant_0(\arbiter|grant[0]~q ),
	.req_and_use_mutex(\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.grant_1(\arbiter|grant[1]~q ),
	.mutex_req(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.grant_7(\arbiter|grant[7]~q ),
	.mutex_req1(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.grant_8(\arbiter|grant[8]~q ),
	.mutex_req2(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.mutex_grant1(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.mutex_grant2(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.mutex_grant3(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.WideNor01(\arbiter|WideNor0~combout ),
	.mgmt_clk_clk(mgmt_clk_clk));

RECONFIGURE_IP_alt_xcvr_reconfig_analog \analog.sc_analog (
	.user_reconfig_readdata_6(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[6]~q ),
	.user_reconfig_readdata_7(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[7]~q ),
	.user_reconfig_readdata_10(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[10]~q ),
	.user_reconfig_readdata_11(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[11]~q ),
	.user_reconfig_readdata_12(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[12]~q ),
	.basic_reconfig_readdata_12(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[12]~q ),
	.user_reconfig_readdata_13(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[13]~q ),
	.basic_reconfig_readdata_13(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[13]~q ),
	.user_reconfig_readdata_14(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[14]~q ),
	.basic_reconfig_readdata_14(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[14]~q ),
	.user_reconfig_readdata_15(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[15]~q ),
	.basic_reconfig_readdata_15(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[15]~q ),
	.user_reconfig_readdata_16(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[16]~q ),
	.basic_reconfig_readdata_16(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[16]~q ),
	.user_reconfig_readdata_17(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[17]~q ),
	.basic_reconfig_readdata_17(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[17]~q ),
	.user_reconfig_readdata_18(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[18]~q ),
	.basic_reconfig_readdata_18(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[18]~q ),
	.user_reconfig_readdata_19(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[19]~q ),
	.basic_reconfig_readdata_19(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[19]~q ),
	.basic_reconfig_readdata_20(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[20]~q ),
	.basic_reconfig_readdata_21(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[21]~q ),
	.basic_reconfig_readdata_22(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[22]~q ),
	.basic_reconfig_readdata_23(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[23]~q ),
	.basic_reconfig_readdata_24(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[24]~q ),
	.basic_reconfig_readdata_25(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[25]~q ),
	.basic_reconfig_readdata_26(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[26]~q ),
	.basic_reconfig_readdata_27(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[27]~q ),
	.basic_reconfig_readdata_28(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[28]~q ),
	.basic_reconfig_readdata_29(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[29]~q ),
	.basic_reconfig_readdata_30(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[30]~q ),
	.basic_reconfig_readdata_31(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[31]~q ),
	.master_writedata_16(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[16]~q ),
	.master_writedata_17(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[17]~q ),
	.master_writedata_18(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[18]~q ),
	.master_writedata_19(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[19]~q ),
	.master_writedata_20(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[20]~q ),
	.master_writedata_21(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[21]~q ),
	.master_writedata_22(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[22]~q ),
	.master_writedata_23(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[23]~q ),
	.master_writedata_24(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[24]~q ),
	.master_writedata_25(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[25]~q ),
	.master_writedata_26(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[26]~q ),
	.master_writedata_27(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[27]~q ),
	.master_writedata_11(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ),
	.master_writedata_28(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[28]~q ),
	.master_writedata_12(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ),
	.master_writedata_29(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[29]~q ),
	.master_writedata_13(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ),
	.master_writedata_30(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[30]~q ),
	.master_writedata_14(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ),
	.master_writedata_31(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[31]~q ),
	.master_writedata_15(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ),
	.rtl(rtl),
	.user_reconfig_readdata_0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[0]~q ),
	.basic_reconfig_readdata_0(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[0]~q ),
	.user_reconfig_readdata_1(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[1]~q ),
	.basic_reconfig_readdata_1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[1]~q ),
	.user_reconfig_readdata_2(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[2]~q ),
	.basic_reconfig_readdata_2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[2]~q ),
	.user_reconfig_readdata_3(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[3]~q ),
	.basic_reconfig_readdata_3(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[3]~q ),
	.user_reconfig_readdata_4(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[4]~q ),
	.basic_reconfig_readdata_4(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[4]~q ),
	.user_reconfig_readdata_5(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[5]~q ),
	.basic_reconfig_readdata_5(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[5]~q ),
	.Equal1(\Equal1~0_combout ),
	.basic_reconfig_readdata_6(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[6]~q ),
	.basic_reconfig_readdata_7(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[7]~q ),
	.basic_reconfig_readdata_8(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[8]~q ),
	.user_reconfig_readdata_8(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[8]~q ),
	.user_reconfig_readdata_9(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_9(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_10(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[10]~q ),
	.basic_reconfig_readdata_11(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[11]~q ),
	.user_reconfig_readdata_20(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[20]~q ),
	.user_reconfig_readdata_21(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[21]~q ),
	.user_reconfig_readdata_22(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[22]~q ),
	.user_reconfig_readdata_23(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[23]~q ),
	.user_reconfig_readdata_24(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[24]~q ),
	.user_reconfig_readdata_25(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[25]~q ),
	.user_reconfig_readdata_26(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[26]~q ),
	.user_reconfig_readdata_27(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[27]~q ),
	.user_reconfig_readdata_28(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[28]~q ),
	.user_reconfig_readdata_29(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[29]~q ),
	.user_reconfig_readdata_30(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[30]~q ),
	.user_reconfig_readdata_31(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[31]~q ),
	.master_write(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_write~q ),
	.grant_1(\arbiter|grant[1]~q ),
	.mutex_req(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.master_address_2(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[2]~q ),
	.mutex_grant(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.master_address_0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ),
	.master_address_1(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[1]~q ),
	.lif_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~1_combout ),
	.master_read(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_read~q ),
	.basic_reconfig_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~0_combout ),
	.basic_reconfig_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~1_combout ),
	.comb(\comb~0_combout ),
	.analog_reconfig_waitrequest(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|wait_gen|wait_req~0_combout ),
	.stateSTATE_IDLE(\analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|inst_analog_ctrlsm|state.STATE_IDLE~q ),
	.ifsel_notdone_resync(\ifsel_notdone_resync~q ),
	.uif_addr_offset_5(uif_addr_offset_5),
	.uif_addr_offset_4(uif_addr_offset_4),
	.uif_addr_offset_0(uif_addr_offset_0),
	.Decoder3(Decoder3),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_1(readdata_for_user_1),
	.Decoder31(Decoder31),
	.Selector2(Selector2),
	.Selector21(Selector21),
	.Decoder32(Decoder32),
	.lpbk_lock(lpbk_lock),
	.analog_offset_0(analog_offset_0),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_9(readdata_for_user_9),
	.rtl1(rtl1),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_13(readdata_for_user_13),
	.rtl2(rtl2),
	.rtl3(rtl3),
	.rtl4(rtl4),
	.rtl5(rtl5),
	.rtl6(rtl6),
	.readdata_for_user_16(readdata_for_user_16),
	.rtl7(rtl7),
	.rtl8(rtl8),
	.WideOr4(WideOr4),
	.WideOr41(WideOr41),
	.analog_length(analog_length),
	.analog_length1(analog_length1),
	.analog_length2(analog_length2),
	.rtl9(rtl9),
	.readdata_for_user_17(readdata_for_user_17),
	.rtl10(rtl10),
	.rtl11(rtl11),
	.user_reconfig_readdata_101(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[10]~7_combout ),
	.rtl12(rtl12),
	.readdata_for_user_18(readdata_for_user_18),
	.rtl13(rtl13),
	.rtl14(rtl14),
	.uif_writedata_4(uif_writedata_4),
	.readdata_for_user_19(readdata_for_user_19),
	.rtl15(rtl15),
	.rtl16(rtl16),
	.LessThan4(LessThan4),
	.readdata_for_user_20(readdata_for_user_20),
	.rtl17(rtl17),
	.rtl18(rtl18),
	.readdata_for_user_21(readdata_for_user_21),
	.rtl19(rtl19),
	.rtl20(rtl20),
	.readdata_for_user_22(readdata_for_user_22),
	.rtl21(rtl21),
	.rtl22(rtl22),
	.readdata_for_user_23(readdata_for_user_23),
	.rtl23(rtl23),
	.readdata_for_user_24(readdata_for_user_24),
	.rtl24(rtl24),
	.readdata_for_user_25(readdata_for_user_25),
	.rtl25(rtl25),
	.readdata_for_user_26(readdata_for_user_26),
	.rtl26(rtl26),
	.readdata_for_user_27(readdata_for_user_27),
	.rtl27(rtl27),
	.readdata_for_user_28(readdata_for_user_28),
	.rtl28(rtl28),
	.readdata_for_user_29(readdata_for_user_29),
	.rtl29(rtl29),
	.readdata_for_user_30(readdata_for_user_30),
	.rtl30(rtl30),
	.readdata_for_user_31(readdata_for_user_31),
	.rtl31(rtl31),
	.rtl32(rtl32),
	.rtl33(rtl33),
	.lif_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~5_combout ),
	.lif_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~6_combout ),
	.Equal8(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|Equal8~0_combout ),
	.basic_reconfig_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~2_combout ),
	.master_writedata_1(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[1]~q ),
	.master_writedata_2(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[2]~q ),
	.master_writedata_0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[0]~q ),
	.master_writedata_3(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[3]~q ),
	.master_writedata_4(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ),
	.master_writedata_5(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ),
	.master_writedata_6(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ),
	.master_writedata_7(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ),
	.master_writedata_8(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ),
	.master_writedata_9(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ),
	.master_writedata_10(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ),
	.uif_mode_0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_mode[0]~0_combout ),
	.Mux0(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux0~0_combout ),
	.Mux3(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux3~0_combout ),
	.WideOr0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|WideOr0~0_combout ),
	.Selector5(Selector5),
	.result_data_0(result_data_0),
	.rtl34(rtl34),
	.rtl35(rtl35),
	.rtl36(rtl36),
	.rtl37(rtl37),
	.rtl38(rtl38),
	.rtl39(rtl39),
	.rtl40(rtl40),
	.rtl41(rtl41),
	.rtl42(rtl42),
	.rtl43(rtl43),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15));

RECONFIGURE_IP_alt_xcvr_reconfig_mif \mif.sc_mif (
	.user_reconfig_readdata_12(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[12]~q ),
	.basic_reconfig_readdata_12(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[12]~q ),
	.user_reconfig_readdata_13(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[13]~q ),
	.basic_reconfig_readdata_13(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[13]~q ),
	.user_reconfig_readdata_14(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[14]~q ),
	.basic_reconfig_readdata_14(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[14]~q ),
	.user_reconfig_readdata_15(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[15]~q ),
	.basic_reconfig_readdata_15(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[15]~q ),
	.user_reconfig_readdata_16(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[16]~q ),
	.basic_reconfig_readdata_16(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[16]~q ),
	.user_reconfig_readdata_17(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[17]~q ),
	.basic_reconfig_readdata_17(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[17]~q ),
	.user_reconfig_readdata_18(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[18]~q ),
	.basic_reconfig_readdata_18(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[18]~q ),
	.user_reconfig_readdata_19(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[19]~q ),
	.basic_reconfig_readdata_19(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[19]~q ),
	.basic_reconfig_readdata_20(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[20]~q ),
	.user_reconfig_readdata_20(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[20]~q ),
	.basic_reconfig_readdata_21(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[21]~q ),
	.user_reconfig_readdata_21(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[21]~q ),
	.basic_reconfig_readdata_22(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[22]~q ),
	.user_reconfig_readdata_22(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[22]~q ),
	.basic_reconfig_readdata_23(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[23]~q ),
	.user_reconfig_readdata_23(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[23]~q ),
	.basic_reconfig_readdata_24(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[24]~q ),
	.user_reconfig_readdata_24(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[24]~q ),
	.basic_reconfig_readdata_25(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[25]~q ),
	.user_reconfig_readdata_25(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[25]~q ),
	.basic_reconfig_readdata_26(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[26]~q ),
	.user_reconfig_readdata_26(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[26]~q ),
	.basic_reconfig_readdata_27(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[27]~q ),
	.user_reconfig_readdata_27(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[27]~q ),
	.basic_reconfig_readdata_28(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[28]~q ),
	.user_reconfig_readdata_28(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[28]~q ),
	.basic_reconfig_readdata_29(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[29]~q ),
	.user_reconfig_readdata_29(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[29]~q ),
	.basic_reconfig_readdata_30(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[30]~q ),
	.user_reconfig_readdata_30(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[30]~q ),
	.basic_reconfig_readdata_31(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[31]~q ),
	.user_reconfig_readdata_31(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[31]~q ),
	.stream_address_0(stream_address_0),
	.stream_address_1(stream_address_1),
	.stream_address_2(stream_address_2),
	.stream_address_3(stream_address_3),
	.stream_address_4(stream_address_4),
	.stream_address_5(stream_address_5),
	.stream_address_6(stream_address_6),
	.stream_address_7(stream_address_7),
	.stream_address_8(stream_address_8),
	.stream_address_9(stream_address_9),
	.stream_address_10(stream_address_10),
	.stream_address_11(stream_address_11),
	.stream_address_12(stream_address_12),
	.stream_address_13(stream_address_13),
	.stream_address_14(stream_address_14),
	.stream_address_15(stream_address_15),
	.stream_address_16(stream_address_16),
	.stream_address_17(stream_address_17),
	.stream_address_18(stream_address_18),
	.stream_address_19(stream_address_19),
	.stream_address_20(stream_address_20),
	.stream_address_21(stream_address_21),
	.stream_address_22(stream_address_22),
	.stream_address_23(stream_address_23),
	.stream_address_24(stream_address_24),
	.stream_address_25(stream_address_25),
	.stream_address_26(stream_address_26),
	.stream_address_27(stream_address_27),
	.stream_address_28(stream_address_28),
	.stream_address_29(stream_address_29),
	.stream_address_30(stream_address_30),
	.stream_address_31(stream_address_31),
	.user_reconfig_readdata_0(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[0]~q ),
	.Equal3(\Equal3~0_combout ),
	.basic_reconfig_readdata_0(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[0]~q ),
	.user_reconfig_readdata_1(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[1]~q ),
	.basic_reconfig_readdata_1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[1]~q ),
	.user_reconfig_readdata_2(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[2]~q ),
	.basic_reconfig_readdata_2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[2]~q ),
	.user_reconfig_readdata_3(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[3]~q ),
	.basic_reconfig_readdata_3(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[3]~q ),
	.user_reconfig_readdata_4(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[4]~q ),
	.basic_reconfig_readdata_4(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[4]~q ),
	.user_reconfig_readdata_5(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[5]~q ),
	.basic_reconfig_readdata_5(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[5]~q ),
	.basic_reconfig_readdata_6(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[6]~q ),
	.user_reconfig_readdata_6(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[6]~q ),
	.basic_reconfig_readdata_7(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[7]~q ),
	.user_reconfig_readdata_7(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[7]~q ),
	.reconfig_mgmt_readdata_8(\reconfig_mgmt_readdata[8]~0_combout ),
	.basic_reconfig_readdata_8(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[8]~q ),
	.user_reconfig_readdata_8(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[8]~q ),
	.user_reconfig_readdata_9(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_9(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_10(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[10]~q ),
	.user_reconfig_readdata_10(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[10]~q ),
	.basic_reconfig_readdata_11(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[11]~q ),
	.user_reconfig_readdata_11(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[11]~q ),
	.master_write(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_write~q ),
	.grant_7(\arbiter|grant[7]~q ),
	.mutex_req(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.mutex_grant(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.master_address_2(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[2]~q ),
	.master_address_0(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ),
	.master_address_1(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[1]~q ),
	.lif_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~1_combout ),
	.master_read(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_read~q ),
	.basic_reconfig_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~0_combout ),
	.basic_reconfig_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~1_combout ),
	.resync_chains0sync_r_1(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ),
	.launch_reg(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|launch_reg~q ),
	.wait_reg(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|wait_reg~q ),
	.stream_read(stream_read),
	.uif_busy(\mif.sc_mif|mif_strm_av|inst_mif_ctrl|uif_busy~q ),
	.pll_mif_busy(\pll.sc_pll|pll_reconfig_av|inst_pll_ctrl|pll_mif_busy~q ),
	.ifsel_notdone_resync(\ifsel_notdone_resync~q ),
	.uif_logical_ch_addr_0(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[0]~q ),
	.comb(\comb~1_combout ),
	.uif_logical_ch_addr_1(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[1]~q ),
	.uif_logical_ch_addr_2(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[2]~q ),
	.uif_logical_ch_addr_3(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[3]~q ),
	.user_reconfig_readdata_101(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[10]~7_combout ),
	.uif_logical_ch_addr_4(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[4]~q ),
	.uif_logical_ch_addr_5(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[5]~q ),
	.uif_logical_ch_addr_6(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[6]~q ),
	.uif_logical_ch_addr_7(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[7]~q ),
	.uif_logical_ch_addr_8(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[8]~q ),
	.uif_logical_ch_addr_9(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[9]~q ),
	.lif_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~5_combout ),
	.lif_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~6_combout ),
	.Equal8(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|Equal8~0_combout ),
	.basic_reconfig_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~2_combout ),
	.master_writedata_1(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[1]~q ),
	.master_writedata_2(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[2]~q ),
	.master_writedata_0(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[0]~q ),
	.master_writedata_3(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[3]~q ),
	.master_writedata_4(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ),
	.master_writedata_5(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ),
	.master_writedata_6(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ),
	.master_writedata_7(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ),
	.master_writedata_8(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ),
	.master_writedata_9(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ),
	.master_writedata_10(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ),
	.master_writedata_11(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ),
	.master_writedata_12(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ),
	.master_writedata_13(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ),
	.master_writedata_14(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ),
	.master_writedata_15(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ),
	.pll_go(\mif.sc_mif|mif_strm_av|inst_mif_avmm|pll_go~q ),
	.uif_mode_0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_mode[0]~0_combout ),
	.Mux0(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux0~0_combout ),
	.Mux3(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux3~0_combout ),
	.WideOr0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|WideOr0~0_combout ),
	.pll_type(\mif.sc_mif|mif_strm_av|inst_mif_avmm|pll_type~q ),
	.mif_rec_addr_7(\mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[7]~q ),
	.mif_rec_addr_5(\mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[5]~q ),
	.mif_rec_addr_6(\mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[6]~q ),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mif_waitrequest(reconfig_mif_waitrequest),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15),
	.reconfig_mif_readdata_15(reconfig_mif_readdata_15),
	.reconfig_mif_readdata_14(reconfig_mif_readdata_14),
	.reconfig_mif_readdata_13(reconfig_mif_readdata_13),
	.reconfig_mif_readdata_12(reconfig_mif_readdata_12),
	.reconfig_mif_readdata_11(reconfig_mif_readdata_11),
	.reconfig_mif_readdata_1(reconfig_mif_readdata_1),
	.reconfig_mif_readdata_0(reconfig_mif_readdata_0),
	.reconfig_mif_readdata_4(reconfig_mif_readdata_4),
	.reconfig_mif_readdata_3(reconfig_mif_readdata_3),
	.reconfig_mif_readdata_2(reconfig_mif_readdata_2),
	.reconfig_mif_readdata_7(reconfig_mif_readdata_7),
	.reconfig_mif_readdata_5(reconfig_mif_readdata_5),
	.reconfig_mif_readdata_6(reconfig_mif_readdata_6),
	.reconfig_mif_readdata_8(reconfig_mif_readdata_8),
	.reconfig_mif_readdata_9(reconfig_mif_readdata_9),
	.reconfig_mif_readdata_10(reconfig_mif_readdata_10));

RECONFIGURE_IP_alt_xcvr_reconfig_direct \direct.sc_direct (
	.Equal2(\Equal2~0_combout ),
	.reg_arb_req1(\direct.sc_direct|reg_arb_req~q ),
	.grant_4(\arbiter|grant[4]~q ),
	.mutex_grant(\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.basic_write(\direct.sc_direct|mutex_inst|master_write~0_combout ),
	.reset(\ifsel_notdone_resync~q ),
	.master_read(\direct.sc_direct|mutex_inst|master_read~combout ),
	.reconfig_mgmt_address_3(reconfig_mgmt_address_3),
	.reconfig_mgmt_address_4(reconfig_mgmt_address_4),
	.reconfig_mgmt_address_5(reconfig_mgmt_address_5),
	.reconfig_mgmt_address_6(reconfig_mgmt_address_6),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0));

RECONFIGURE_IP_alt_xcvr_reconfig_cal_seq cal_seq(
	.reconfig_busy1(reconfig_busy),
	.offset_cancellation_done(offset_cancellation_done),
	.tx_cal_busy1(tx_cal_busy),
	.rx_cal_busy1(rx_cal_busy),
	.uif_busy(\mif.sc_mif|mif_strm_av|inst_mif_ctrl|uif_busy~q ),
	.pll_mif_busy(\pll.sc_pll|pll_reconfig_av|inst_pll_ctrl|pll_mif_busy~q ),
	.stateSTATE_IDLE(\analog.sc_analog|reconfig_analog_cv|inst_analog_datactrl|inst_analog_ctrlsm|state.STATE_IDLE~q ),
	.ifsel_notdone_resync(\ifsel_notdone_resync~q ),
	.mgmt_clk_clk(mgmt_clk_clk));

RECONFIGURE_IP_alt_xcvr_reconfig_pll \pll.sc_pll (
	.user_reconfig_readdata_10(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[10]~q ),
	.user_reconfig_readdata_11(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[11]~q ),
	.user_reconfig_readdata_12(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[12]~q ),
	.basic_reconfig_readdata_12(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[12]~q ),
	.user_reconfig_readdata_13(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[13]~q ),
	.basic_reconfig_readdata_13(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[13]~q ),
	.user_reconfig_readdata_14(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[14]~q ),
	.basic_reconfig_readdata_14(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[14]~q ),
	.user_reconfig_readdata_15(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[15]~q ),
	.basic_reconfig_readdata_15(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[15]~q ),
	.user_reconfig_readdata_16(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[16]~q ),
	.basic_reconfig_readdata_16(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[16]~q ),
	.user_reconfig_readdata_17(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[17]~q ),
	.basic_reconfig_readdata_17(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[17]~q ),
	.user_reconfig_readdata_18(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[18]~q ),
	.basic_reconfig_readdata_18(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[18]~q ),
	.user_reconfig_readdata_19(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[19]~q ),
	.basic_reconfig_readdata_19(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[19]~q ),
	.basic_reconfig_readdata_20(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[20]~q ),
	.user_reconfig_readdata_20(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[20]~q ),
	.basic_reconfig_readdata_21(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[21]~q ),
	.user_reconfig_readdata_21(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[21]~q ),
	.basic_reconfig_readdata_22(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[22]~q ),
	.user_reconfig_readdata_22(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[22]~q ),
	.basic_reconfig_readdata_23(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[23]~q ),
	.user_reconfig_readdata_23(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[23]~q ),
	.basic_reconfig_readdata_24(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[24]~q ),
	.user_reconfig_readdata_24(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[24]~q ),
	.basic_reconfig_readdata_25(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[25]~q ),
	.basic_reconfig_readdata_26(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[26]~q ),
	.basic_reconfig_readdata_27(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[27]~q ),
	.basic_reconfig_readdata_28(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[28]~q ),
	.basic_reconfig_readdata_29(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[29]~q ),
	.basic_reconfig_readdata_30(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[30]~q ),
	.basic_reconfig_readdata_31(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[31]~q ),
	.user_reconfig_readdata_0(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[0]~q ),
	.Equal4(\Equal4~0_combout ),
	.basic_reconfig_readdata_0(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[0]~q ),
	.user_reconfig_readdata_1(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[1]~q ),
	.basic_reconfig_readdata_1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[1]~q ),
	.user_reconfig_readdata_2(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[2]~q ),
	.basic_reconfig_readdata_2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[2]~q ),
	.user_reconfig_readdata_3(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[3]~q ),
	.basic_reconfig_readdata_3(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[3]~q ),
	.user_reconfig_readdata_4(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[4]~q ),
	.basic_reconfig_readdata_4(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[4]~q ),
	.user_reconfig_readdata_5(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[5]~q ),
	.basic_reconfig_readdata_5(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[5]~q ),
	.basic_reconfig_readdata_6(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[6]~q ),
	.user_reconfig_readdata_6(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[6]~q ),
	.basic_reconfig_readdata_7(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[7]~q ),
	.user_reconfig_readdata_7(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[7]~q ),
	.user_reconfig_readdata_8(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[8]~q ),
	.basic_reconfig_readdata_8(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[8]~q ),
	.user_reconfig_readdata_9(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_9(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_10(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[10]~q ),
	.basic_reconfig_readdata_11(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[11]~q ),
	.user_reconfig_readdata_25(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[25]~q ),
	.user_reconfig_readdata_26(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[26]~q ),
	.user_reconfig_readdata_27(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[27]~q ),
	.user_reconfig_readdata_28(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[28]~q ),
	.user_reconfig_readdata_29(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[29]~q ),
	.user_reconfig_readdata_30(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[30]~q ),
	.user_reconfig_readdata_31(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[31]~q ),
	.master_write(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_write~q ),
	.grant_8(\arbiter|grant[8]~q ),
	.mutex_req(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.master_address_2(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_address[2]~combout ),
	.master_address_0(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ),
	.master_address_1(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_address[1]~combout ),
	.lif_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~1_combout ),
	.master_read(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_read~q ),
	.basic_reconfig_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~0_combout ),
	.basic_reconfig_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~1_combout ),
	.resync_chains0sync_r_1(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ),
	.launch_reg(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|launch_reg~q ),
	.wait_reg(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|wait_reg~q ),
	.pll_mif_busy(\pll.sc_pll|pll_reconfig_av|inst_pll_ctrl|pll_mif_busy~q ),
	.ifsel_notdone_resync(\ifsel_notdone_resync~q ),
	.uif_logical_ch_addr_0(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[0]~q ),
	.comb(\comb~2_combout ),
	.uif_logical_ch_addr_1(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[1]~q ),
	.uif_logical_ch_addr_2(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[2]~q ),
	.uif_logical_ch_addr_3(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[3]~q ),
	.user_reconfig_readdata_101(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[10]~7_combout ),
	.uif_logical_ch_addr_4(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[4]~q ),
	.uif_logical_ch_addr_5(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[5]~q ),
	.uif_logical_ch_addr_6(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[6]~q ),
	.uif_logical_ch_addr_7(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[7]~q ),
	.uif_logical_ch_addr_8(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[8]~q ),
	.uif_logical_ch_addr_9(\mif.sc_mif|mif_strm_av|inst_xreconf_uif|uif_logical_ch_addr[9]~q ),
	.mutex_grant(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.lif_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~5_combout ),
	.lif_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~6_combout ),
	.Equal8(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|Equal8~0_combout ),
	.basic_reconfig_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~2_combout ),
	.master_writedata_1(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[1]~combout ),
	.master_writedata_2(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[2]~combout ),
	.master_writedata_0(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[0]~combout ),
	.master_writedata_3(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[3]~combout ),
	.master_writedata_4(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ),
	.master_writedata_5(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ),
	.master_writedata_6(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ),
	.master_writedata_7(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ),
	.master_writedata_8(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ),
	.master_writedata_9(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ),
	.master_writedata_10(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ),
	.master_writedata_11(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ),
	.master_writedata_12(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ),
	.master_writedata_13(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ),
	.master_writedata_14(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ),
	.master_writedata_15(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ),
	.pll_go(\mif.sc_mif|mif_strm_av|inst_mif_avmm|pll_go~q ),
	.uif_mode_0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|uif_mode[0]~0_combout ),
	.Mux0(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux0~0_combout ),
	.Mux3(\pll.sc_pll|pll_reconfig_av|inst_pll_uif|Mux3~0_combout ),
	.WideOr0(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|WideOr0~0_combout ),
	.pll_type(\mif.sc_mif|mif_strm_av|inst_mif_avmm|pll_type~q ),
	.mif_rec_addr_7(\mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[7]~q ),
	.mif_rec_addr_5(\mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[5]~q ),
	.mif_rec_addr_6(\mif.sc_mif|mif_strm_av|inst_mif_avmm|mif_rec_addr[6]~q ),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15));

RECONFIGURE_IP_alt_xcvr_reconfig_basic basic(
	.basic_reconfig_readdata_12(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[12]~q ),
	.basic_reconfig_readdata_13(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[13]~q ),
	.basic_reconfig_readdata_14(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[14]~q ),
	.basic_reconfig_readdata_15(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[15]~q ),
	.basic_reconfig_readdata_16(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[16]~q ),
	.basic_reconfig_readdata_17(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[17]~q ),
	.basic_reconfig_readdata_18(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[18]~q ),
	.basic_reconfig_readdata_19(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[19]~q ),
	.basic_reconfig_readdata_20(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[20]~q ),
	.basic_reconfig_readdata_21(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[21]~q ),
	.basic_reconfig_readdata_22(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[22]~q ),
	.basic_reconfig_readdata_23(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[23]~q ),
	.basic_reconfig_readdata_24(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[24]~q ),
	.basic_reconfig_readdata_25(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[25]~q ),
	.basic_reconfig_readdata_26(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[26]~q ),
	.basic_reconfig_readdata_27(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[27]~q ),
	.basic_reconfig_readdata_28(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[28]~q ),
	.basic_reconfig_readdata_29(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[29]~q ),
	.basic_reconfig_readdata_30(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[30]~q ),
	.basic_reconfig_readdata_31(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[31]~q ),
	.master_writedata_16(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[16]~q ),
	.master_writedata_17(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[17]~q ),
	.master_writedata_18(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[18]~q ),
	.master_writedata_19(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[19]~q ),
	.master_writedata_20(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[20]~q ),
	.master_writedata_21(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[21]~q ),
	.master_writedata_22(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[22]~q ),
	.master_writedata_23(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[23]~q ),
	.master_writedata_24(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[24]~q ),
	.master_writedata_25(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[25]~q ),
	.master_writedata_26(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[26]~q ),
	.master_writedata_27(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[27]~q ),
	.master_writedata_28(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[28]~q ),
	.master_writedata_12(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ),
	.master_writedata_29(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[29]~q ),
	.master_writedata_13(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ),
	.master_writedata_30(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[30]~q ),
	.master_writedata_14(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ),
	.master_writedata_31(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[31]~q ),
	.master_writedata_15(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ),
	.basic_reconfig_readdata_0(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[0]~q ),
	.basic_reconfig_readdata_1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[1]~q ),
	.basic_reconfig_readdata_2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[2]~q ),
	.basic_reconfig_readdata_3(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[3]~q ),
	.basic_reconfig_readdata_4(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[4]~q ),
	.basic_reconfig_readdata_5(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[5]~q ),
	.Equal2(\Equal2~0_combout ),
	.basic_reconfig_readdata_6(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[6]~q ),
	.basic_reconfig_readdata_7(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[7]~q ),
	.basic_reconfig_readdata_8(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[8]~q ),
	.basic_reconfig_readdata_9(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[9]~q ),
	.basic_reconfig_readdata_10(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[10]~q ),
	.basic_reconfig_readdata_11(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[11]~q ),
	.mutex_grant(\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.master_write(\direct.sc_direct|mutex_inst|master_write~0_combout ),
	.wbasic_write_8(\wbasic_write[8]~0_combout ),
	.wbasic_write_81(\wbasic_write[8]~1_combout ),
	.wbasic_write_82(\wbasic_write[8]~2_combout ),
	.mutex_grant1(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.wbasic_address_2_8(\wbasic_address[8][2]~combout ),
	.mutex_grant2(\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.wbasic_address_0_8(\wbasic_address[8][0]~3_combout ),
	.wbasic_address_1_8(\wbasic_address[8][1]~combout ),
	.lif_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~1_combout ),
	.wbasic_read_8(\wbasic_read[8]~0_combout ),
	.wbasic_read_81(\wbasic_read[8]~1_combout ),
	.basic_reconfig_waitrequest(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~0_combout ),
	.basic_reconfig_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~1_combout ),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.native_reconfig_writedata_0(native_reconfig_writedata_0),
	.native_reconfig_writedata_1(native_reconfig_writedata_1),
	.native_reconfig_writedata_2(native_reconfig_writedata_2),
	.native_reconfig_writedata_3(native_reconfig_writedata_3),
	.native_reconfig_writedata_4(native_reconfig_writedata_4),
	.native_reconfig_writedata_5(native_reconfig_writedata_5),
	.native_reconfig_writedata_6(native_reconfig_writedata_6),
	.native_reconfig_writedata_7(native_reconfig_writedata_7),
	.native_reconfig_writedata_8(native_reconfig_writedata_8),
	.native_reconfig_writedata_9(native_reconfig_writedata_9),
	.native_reconfig_writedata_10(native_reconfig_writedata_10),
	.native_reconfig_writedata_11(native_reconfig_writedata_11),
	.native_reconfig_writedata_12(native_reconfig_writedata_12),
	.native_reconfig_writedata_13(native_reconfig_writedata_13),
	.native_reconfig_writedata_14(native_reconfig_writedata_14),
	.native_reconfig_writedata_15(native_reconfig_writedata_15),
	.native_reconfig_write_0(native_reconfig_write_0),
	.native_reconfig_read_0(native_reconfig_read_0),
	.native_reconfig_address_0(native_reconfig_address_0),
	.native_reconfig_address_1(native_reconfig_address_1),
	.native_reconfig_address_2(native_reconfig_address_2),
	.native_reconfig_address_3(native_reconfig_address_3),
	.native_reconfig_address_4(native_reconfig_address_4),
	.native_reconfig_address_5(native_reconfig_address_5),
	.native_reconfig_address_6(native_reconfig_address_6),
	.native_reconfig_address_7(native_reconfig_address_7),
	.native_reconfig_address_8(native_reconfig_address_8),
	.native_reconfig_address_9(native_reconfig_address_9),
	.native_reconfig_address_10(native_reconfig_address_10),
	.native_reconfig_address_11(native_reconfig_address_11),
	.pif_testbus_sel_0(pif_testbus_sel_0),
	.pif_testbus_sel_1(pif_testbus_sel_1),
	.pif_testbus_sel_2(pif_testbus_sel_2),
	.pif_testbus_sel_3(pif_testbus_sel_3),
	.pif_interface_sel(pif_interface_sel),
	.pif_ser_shift_load(pif_ser_shift_load),
	.native_reconfig_writedata_16(native_reconfig_writedata_16),
	.native_reconfig_writedata_17(native_reconfig_writedata_17),
	.native_reconfig_writedata_18(native_reconfig_writedata_18),
	.native_reconfig_writedata_19(native_reconfig_writedata_19),
	.native_reconfig_writedata_20(native_reconfig_writedata_20),
	.native_reconfig_writedata_21(native_reconfig_writedata_21),
	.native_reconfig_writedata_22(native_reconfig_writedata_22),
	.native_reconfig_writedata_23(native_reconfig_writedata_23),
	.native_reconfig_writedata_24(native_reconfig_writedata_24),
	.native_reconfig_writedata_25(native_reconfig_writedata_25),
	.native_reconfig_writedata_26(native_reconfig_writedata_26),
	.native_reconfig_writedata_27(native_reconfig_writedata_27),
	.native_reconfig_writedata_28(native_reconfig_writedata_28),
	.native_reconfig_writedata_29(native_reconfig_writedata_29),
	.native_reconfig_writedata_30(native_reconfig_writedata_30),
	.native_reconfig_writedata_31(native_reconfig_writedata_31),
	.native_reconfig_write_1(native_reconfig_write_1),
	.native_reconfig_read_1(native_reconfig_read_1),
	.native_reconfig_address_12(native_reconfig_address_12),
	.native_reconfig_address_13(native_reconfig_address_13),
	.native_reconfig_address_14(native_reconfig_address_14),
	.native_reconfig_address_15(native_reconfig_address_15),
	.native_reconfig_address_16(native_reconfig_address_16),
	.native_reconfig_address_17(native_reconfig_address_17),
	.native_reconfig_address_18(native_reconfig_address_18),
	.native_reconfig_address_19(native_reconfig_address_19),
	.native_reconfig_address_20(native_reconfig_address_20),
	.native_reconfig_address_21(native_reconfig_address_21),
	.native_reconfig_address_22(native_reconfig_address_22),
	.native_reconfig_address_23(native_reconfig_address_23),
	.pif_testbus_sel_12(pif_testbus_sel_12),
	.pif_testbus_sel_13(pif_testbus_sel_13),
	.pif_testbus_sel_14(pif_testbus_sel_14),
	.pif_testbus_sel_15(pif_testbus_sel_15),
	.mutex_grant3(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.mutex_grant4(\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.lif_waitrequest1(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~5_combout ),
	.master_read(\direct.sc_direct|mutex_inst|master_read~combout ),
	.wbasic_read_82(\wbasic_read[8]~2_combout ),
	.lif_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~6_combout ),
	.basic_reconfig_waitrequest2(\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~2_combout ),
	.wbasic_writedata_1_8(\wbasic_writedata[8][1]~combout ),
	.wbasic_writedata_2_8(\wbasic_writedata[8][2]~combout ),
	.wbasic_writedata_0_8(\wbasic_writedata[8][0]~combout ),
	.wbasic_writedata_3_8(\wbasic_writedata[8][3]~combout ),
	.wbasic_writedata_4_8(\wbasic_writedata[8][4]~combout ),
	.wbasic_writedata_5_8(\wbasic_writedata[8][5]~combout ),
	.wbasic_writedata_6_8(\wbasic_writedata[8][6]~combout ),
	.wbasic_writedata_7_8(\wbasic_writedata[8][7]~combout ),
	.wbasic_writedata_8_8(\wbasic_writedata[8][8]~combout ),
	.wbasic_writedata_9_8(\wbasic_writedata[8][9]~combout ),
	.wbasic_writedata_10_8(\wbasic_writedata[8][10]~combout ),
	.wbasic_writedata_11_8(\wbasic_writedata[8][11]~combout ),
	.master_writedata_121(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ),
	.master_write_data_12(\offset.sc_offset|offset_cancellation_av|master_write_data[12]~q ),
	.master_writedata_122(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[12]~q ),
	.master_writedata_131(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ),
	.master_write_data_13(\offset.sc_offset|offset_cancellation_av|master_write_data[13]~q ),
	.master_writedata_132(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[13]~q ),
	.master_writedata_141(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ),
	.master_write_data_14(\offset.sc_offset|offset_cancellation_av|master_write_data[14]~q ),
	.master_writedata_142(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[14]~q ),
	.master_writedata_151(\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ),
	.master_write_data_15(\offset.sc_offset|offset_cancellation_av|master_write_data[15]~q ),
	.master_writedata_152(\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[15]~q ),
	.LessThan0(\basic|a5|LessThan0~0_combout ),
	.wbasic_write_83(\wbasic_write[8]~combout ),
	.lif_is_active(\lif_is_active~combout ),
	.out_narrow_0(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[0]~combout ),
	.out_narrow_1(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[1]~combout ),
	.out_narrow_2(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[2]~combout ),
	.out_narrow_3(\basic|a5|lif[0].logical_if|pif_tbus_mux|out_narrow[3]~combout ),
	.GND_port(GND_port),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_from_xcvr_0(reconfig_from_xcvr_0),
	.reconfig_from_xcvr_46(reconfig_from_xcvr_46),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_from_xcvr_1(reconfig_from_xcvr_1),
	.reconfig_from_xcvr_47(reconfig_from_xcvr_47),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_from_xcvr_2(reconfig_from_xcvr_2),
	.reconfig_from_xcvr_48(reconfig_from_xcvr_48),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_from_xcvr_3(reconfig_from_xcvr_3),
	.reconfig_from_xcvr_49(reconfig_from_xcvr_49),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_from_xcvr_4(reconfig_from_xcvr_4),
	.reconfig_from_xcvr_50(reconfig_from_xcvr_50),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_from_xcvr_5(reconfig_from_xcvr_5),
	.reconfig_from_xcvr_51(reconfig_from_xcvr_51),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_from_xcvr_6(reconfig_from_xcvr_6),
	.reconfig_from_xcvr_52(reconfig_from_xcvr_52),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_from_xcvr_7(reconfig_from_xcvr_7),
	.reconfig_from_xcvr_53(reconfig_from_xcvr_53),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_from_xcvr_8(reconfig_from_xcvr_8),
	.reconfig_from_xcvr_54(reconfig_from_xcvr_54),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_from_xcvr_9(reconfig_from_xcvr_9),
	.reconfig_from_xcvr_55(reconfig_from_xcvr_55),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_from_xcvr_10(reconfig_from_xcvr_10),
	.reconfig_from_xcvr_56(reconfig_from_xcvr_56),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_from_xcvr_11(reconfig_from_xcvr_11),
	.reconfig_from_xcvr_57(reconfig_from_xcvr_57),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_from_xcvr_12(reconfig_from_xcvr_12),
	.reconfig_from_xcvr_58(reconfig_from_xcvr_58),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_from_xcvr_13(reconfig_from_xcvr_13),
	.reconfig_from_xcvr_59(reconfig_from_xcvr_59),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_from_xcvr_14(reconfig_from_xcvr_14),
	.reconfig_from_xcvr_60(reconfig_from_xcvr_60),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15),
	.reconfig_from_xcvr_15(reconfig_from_xcvr_15),
	.reconfig_from_xcvr_61(reconfig_from_xcvr_61),
	.reconfig_from_xcvr_24(reconfig_from_xcvr_24),
	.reconfig_from_xcvr_70(reconfig_from_xcvr_70),
	.reconfig_from_xcvr_16(reconfig_from_xcvr_16),
	.reconfig_from_xcvr_62(reconfig_from_xcvr_62),
	.reconfig_from_xcvr_32(reconfig_from_xcvr_32),
	.reconfig_from_xcvr_78(reconfig_from_xcvr_78),
	.reconfig_from_xcvr_25(reconfig_from_xcvr_25),
	.reconfig_from_xcvr_71(reconfig_from_xcvr_71),
	.reconfig_from_xcvr_17(reconfig_from_xcvr_17),
	.reconfig_from_xcvr_63(reconfig_from_xcvr_63),
	.reconfig_from_xcvr_33(reconfig_from_xcvr_33),
	.reconfig_from_xcvr_79(reconfig_from_xcvr_79),
	.reconfig_from_xcvr_26(reconfig_from_xcvr_26),
	.reconfig_from_xcvr_72(reconfig_from_xcvr_72),
	.reconfig_from_xcvr_18(reconfig_from_xcvr_18),
	.reconfig_from_xcvr_64(reconfig_from_xcvr_64),
	.reconfig_from_xcvr_34(reconfig_from_xcvr_34),
	.reconfig_from_xcvr_80(reconfig_from_xcvr_80),
	.reconfig_from_xcvr_27(reconfig_from_xcvr_27),
	.reconfig_from_xcvr_73(reconfig_from_xcvr_73),
	.reconfig_from_xcvr_19(reconfig_from_xcvr_19),
	.reconfig_from_xcvr_65(reconfig_from_xcvr_65),
	.reconfig_from_xcvr_35(reconfig_from_xcvr_35),
	.reconfig_from_xcvr_81(reconfig_from_xcvr_81));

cyclonev_lcell_comb \wbasic_write[8]~0 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|master_write~q ),
	.datab(!\arbiter|grant[0]~q ),
	.datac(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_write~q ),
	.datae(!\arbiter|grant[1]~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_write[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_write[8]~0 .extended_lut = "off";
defparam \wbasic_write[8]~0 .lut_mask = 64'h01010101010101FF;
defparam \wbasic_write[8]~0 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_write[8]~1 (
	.dataa(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_write~q ),
	.datab(!\arbiter|grant[7]~q ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_write~q ),
	.datae(!\arbiter|grant[8]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_write[8]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_write[8]~1 .extended_lut = "off";
defparam \wbasic_write[8]~1 .lut_mask = 64'h01010101010101FF;
defparam \wbasic_write[8]~1 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_write[8]~2 (
	.dataa(!\wbasic_write[8]~0_combout ),
	.datab(!\wbasic_write[8]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_write[8]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_write[8]~2 .extended_lut = "off";
defparam \wbasic_write[8]~2 .lut_mask = 64'h8888888888888888;
defparam \wbasic_write[8]~2 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_address[8][2]~0 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\arbiter|grant[1]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|master_address[2]~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_address[8][2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_address[8][2]~0 .extended_lut = "off";
defparam \wbasic_address[8][2]~0 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_address[8][2]~0 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_address[8][2] (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[2]~q ),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_address[2]~combout ),
	.dataf(!\wbasic_address[8][2]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_address[8][2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_address[8][2] .extended_lut = "off";
defparam \wbasic_address[8][2] .lut_mask = 64'hEEE0000000000000;
defparam \wbasic_address[8][2] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_address[8][0]~1 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_address[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_address[8][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_address[8][0]~1 .extended_lut = "off";
defparam \wbasic_address[8][0]~1 .lut_mask = 64'h0101010101010101;
defparam \wbasic_address[8][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_address[8][0]~2 (
	.dataa(!\arbiter|grant[7]~q ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datac(!\arbiter|grant[8]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_address[8][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_address[8][0]~2 .extended_lut = "off";
defparam \wbasic_address[8][0]~2 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_address[8][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_address[8][0]~3 (
	.dataa(!reconfig_mgmt_address_0),
	.datab(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[0]~q ),
	.datae(!\wbasic_address[8][0]~1_combout ),
	.dataf(!\wbasic_address[8][0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_address[8][0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_address[8][0]~3 .extended_lut = "off";
defparam \wbasic_address[8][0]~3 .lut_mask = 64'hEEE0000000000000;
defparam \wbasic_address[8][0]~3 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_address[8][1]~4 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\arbiter|grant[1]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|master_address[1]~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_address[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_address[8][1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_address[8][1]~4 .extended_lut = "off";
defparam \wbasic_address[8][1]~4 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_address[8][1]~4 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_address[8][1] (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_address[1]~q ),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_address[1]~combout ),
	.dataf(!\wbasic_address[8][1]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_address[8][1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_address[8][1] .extended_lut = "off";
defparam \wbasic_address[8][1] .lut_mask = 64'hEEE0000000000000;
defparam \wbasic_address[8][1] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_read[8]~0 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\arbiter|grant[1]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|master_read~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_read~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_read[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_read[8]~0 .extended_lut = "off";
defparam \wbasic_read[8]~0 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_read[8]~0 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_read[8]~1 (
	.dataa(!\arbiter|grant[7]~q ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datac(!\arbiter|grant[8]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_read~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_read~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_read[8]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_read[8]~1 .extended_lut = "off";
defparam \wbasic_read[8]~1 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_read[8]~1 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!reconfig_mgmt_read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h0000400000004000;
defparam \comb~0 .shared_arith = "off";

dffeas ifsel_notdone_resync(
	.clk(mgmt_clk_clk),
	.d(\basic|a5|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(resync_chains0sync_r_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ifsel_notdone_resync~q ),
	.prn(vcc));
defparam ifsel_notdone_resync.is_wysiwyg = "true";
defparam ifsel_notdone_resync.power_up = "low";

cyclonev_lcell_comb \comb~1 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!reconfig_mgmt_read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~1 .extended_lut = "off";
defparam \comb~1 .lut_mask = 64'h0000010000000100;
defparam \comb~1 .shared_arith = "off";

cyclonev_lcell_comb \comb~2 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!reconfig_mgmt_read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~2 .extended_lut = "off";
defparam \comb~2 .lut_mask = 64'h0000008000000080;
defparam \comb~2 .shared_arith = "off";

cyclonev_lcell_comb \comb~3 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!reconfig_mgmt_read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~3 .extended_lut = "off";
defparam \comb~3 .lut_mask = 64'h0000800000008000;
defparam \comb~3 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_read[8]~2 (
	.dataa(!\wbasic_read[8]~0_combout ),
	.datab(!\wbasic_read[8]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_read[8]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_read[8]~2 .extended_lut = "off";
defparam \wbasic_read[8]~2 .lut_mask = 64'h8888888888888888;
defparam \wbasic_read[8]~2 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][1]~0 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\arbiter|grant[1]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|master_write_data[1]~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][1]~0 .extended_lut = "off";
defparam \wbasic_writedata[8][1]~0 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_writedata[8][1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][1] (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_1),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[1]~q ),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[1]~combout ),
	.dataf(!\wbasic_writedata[8][1]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][1] .extended_lut = "off";
defparam \wbasic_writedata[8][1] .lut_mask = 64'h0537FFFFFFFFFFFF;
defparam \wbasic_writedata[8][1] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][2]~1 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\arbiter|grant[1]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|master_write_data[2]~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][2]~1 .extended_lut = "off";
defparam \wbasic_writedata[8][2]~1 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_writedata[8][2]~1 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][2] (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_2),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[2]~q ),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[2]~combout ),
	.dataf(!\wbasic_writedata[8][2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][2] .extended_lut = "off";
defparam \wbasic_writedata[8][2] .lut_mask = 64'h0537FFFFFFFFFFFF;
defparam \wbasic_writedata[8][2] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][0]~2 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\arbiter|grant[1]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|master_write_data[0]~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][0]~2 .extended_lut = "off";
defparam \wbasic_writedata[8][0]~2 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_writedata[8][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][0] (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_0),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[0]~q ),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[0]~combout ),
	.dataf(!\wbasic_writedata[8][0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][0] .extended_lut = "off";
defparam \wbasic_writedata[8][0] .lut_mask = 64'h0537FFFFFFFFFFFF;
defparam \wbasic_writedata[8][0] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][3]~3 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\offset.sc_offset|offset_cancellation_av|req_and_use_mutex~q ),
	.datac(!\arbiter|grant[1]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|mutex_req~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|master_write_data[3]~q ),
	.dataf(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][3]~3 .extended_lut = "off";
defparam \wbasic_writedata[8][3]~3 .lut_mask = 64'h00001111000F111F;
defparam \wbasic_writedata[8][3]~3 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][3] (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_3),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[3]~q ),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|master_writedata[3]~combout ),
	.dataf(!\wbasic_writedata[8][3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][3] .extended_lut = "off";
defparam \wbasic_writedata[8][3] .lut_mask = 64'h0537FFFFFFFFFFFF;
defparam \wbasic_writedata[8][3] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][4]~4 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[4]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][4]~4 .extended_lut = "off";
defparam \wbasic_writedata[8][4]~4 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][4]~4 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][4]~5 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_4),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][4]~5 .extended_lut = "off";
defparam \wbasic_writedata[8][4]~5 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][4]~5 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][4] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[4]~q ),
	.datac(!\wbasic_writedata[8][4]~4_combout ),
	.datad(!\wbasic_writedata[8][4]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][4] .extended_lut = "off";
defparam \wbasic_writedata[8][4] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \wbasic_writedata[8][4] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][5]~6 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[5]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][5]~6 .extended_lut = "off";
defparam \wbasic_writedata[8][5]~6 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][5]~6 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][5]~7 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_5),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][5]~7 .extended_lut = "off";
defparam \wbasic_writedata[8][5]~7 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][5]~7 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][5] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[5]~q ),
	.datac(!\wbasic_writedata[8][5]~6_combout ),
	.datad(!\wbasic_writedata[8][5]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][5] .extended_lut = "off";
defparam \wbasic_writedata[8][5] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \wbasic_writedata[8][5] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][6]~8 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[6]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][6]~8 .extended_lut = "off";
defparam \wbasic_writedata[8][6]~8 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][6]~8 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][6]~9 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_6),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][6]~9 .extended_lut = "off";
defparam \wbasic_writedata[8][6]~9 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][6]~9 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][6] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[6]~q ),
	.datac(!\wbasic_writedata[8][6]~8_combout ),
	.datad(!\wbasic_writedata[8][6]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][6] .extended_lut = "off";
defparam \wbasic_writedata[8][6] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \wbasic_writedata[8][6] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][7]~10 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[7]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][7]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][7]~10 .extended_lut = "off";
defparam \wbasic_writedata[8][7]~10 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][7]~10 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][7]~11 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_7),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][7]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][7]~11 .extended_lut = "off";
defparam \wbasic_writedata[8][7]~11 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][7]~11 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][7] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[7]~q ),
	.datac(!\wbasic_writedata[8][7]~10_combout ),
	.datad(!\wbasic_writedata[8][7]~11_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][7] .extended_lut = "off";
defparam \wbasic_writedata[8][7] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \wbasic_writedata[8][7] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][8]~12 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[8]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][8]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][8]~12 .extended_lut = "off";
defparam \wbasic_writedata[8][8]~12 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][8]~12 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][8]~13 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_8),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][8]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][8]~13 .extended_lut = "off";
defparam \wbasic_writedata[8][8]~13 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][8]~13 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][8] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[8]~q ),
	.datac(!\wbasic_writedata[8][8]~12_combout ),
	.datad(!\wbasic_writedata[8][8]~13_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][8] .extended_lut = "off";
defparam \wbasic_writedata[8][8] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \wbasic_writedata[8][8] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][9]~14 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[9]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][9]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][9]~14 .extended_lut = "off";
defparam \wbasic_writedata[8][9]~14 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][9]~14 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][9]~15 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_9),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][9]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][9]~15 .extended_lut = "off";
defparam \wbasic_writedata[8][9]~15 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][9]~15 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][9] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[9]~q ),
	.datac(!\wbasic_writedata[8][9]~14_combout ),
	.datad(!\wbasic_writedata[8][9]~15_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][9] .extended_lut = "off";
defparam \wbasic_writedata[8][9] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \wbasic_writedata[8][9] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][10]~16 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[10]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][10]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][10]~16 .extended_lut = "off";
defparam \wbasic_writedata[8][10]~16 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][10]~16 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][10]~17 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_10),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][10]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][10]~17 .extended_lut = "off";
defparam \wbasic_writedata[8][10]~17 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][10]~17 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][10] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[10]~q ),
	.datac(!\wbasic_writedata[8][10]~16_combout ),
	.datad(!\wbasic_writedata[8][10]~17_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][10] .extended_lut = "off";
defparam \wbasic_writedata[8][10] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \wbasic_writedata[8][10] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][11]~18 (
	.dataa(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datab(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_writedata_11),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][11]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][11]~18 .extended_lut = "off";
defparam \wbasic_writedata[8][11]~18 .lut_mask = 64'h0537053705370537;
defparam \wbasic_writedata[8][11]~18 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][11]~19 (
	.dataa(!\offset.sc_offset|offset_cancellation_av|mutex_inst|mutex_grant~0_combout ),
	.datab(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datac(!\offset.sc_offset|offset_cancellation_av|master_write_data[11]~q ),
	.datad(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ),
	.datae(!\wbasic_writedata[8][11]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][11]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][11]~19 .extended_lut = "off";
defparam \wbasic_writedata[8][11]~19 .lut_mask = 64'hFAC80000FAC80000;
defparam \wbasic_writedata[8][11]~19 .shared_arith = "off";

cyclonev_lcell_comb \wbasic_writedata[8][11] (
	.dataa(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|mutex_inst|mutex_grant~combout ),
	.datab(!\pll.sc_pll|pll_reconfig_av|inst_xreconf_cif|inst_basic_acq|master_writedata[11]~q ),
	.datac(!\wbasic_writedata[8][11]~19_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_writedata[8][11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_writedata[8][11] .extended_lut = "off";
defparam \wbasic_writedata[8][11] .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \wbasic_writedata[8][11] .shared_arith = "off";

cyclonev_lcell_comb \wbasic_write[8] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\direct.sc_direct|mutex_inst|mutex_grant~combout ),
	.datac(!reconfig_mgmt_write),
	.datad(!\wbasic_write[8]~0_combout ),
	.datae(!\wbasic_write[8]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wbasic_write[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wbasic_write[8] .extended_lut = "off";
defparam \wbasic_write[8] .lut_mask = 64'hFE000000FE000000;
defparam \wbasic_write[8] .shared_arith = "off";

dffeas \reg_grant_last[4] (
	.clk(mgmt_clk_clk),
	.d(\arbiter|grant[4]~q ),
	.asdata(vcc),
	.clrn(resync_chains0sync_r_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reg_grant_last[4]~q ),
	.prn(vcc));
defparam \reg_grant_last[4] .is_wysiwyg = "true";
defparam \reg_grant_last[4] .power_up = "low";

dffeas \reg_grant_last[7] (
	.clk(mgmt_clk_clk),
	.d(\arbiter|grant[7]~q ),
	.asdata(vcc),
	.clrn(resync_chains0sync_r_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reg_grant_last[7]~q ),
	.prn(vcc));
defparam \reg_grant_last[7] .is_wysiwyg = "true";
defparam \reg_grant_last[7] .power_up = "low";

dffeas \reg_grant_last[8] (
	.clk(mgmt_clk_clk),
	.d(\arbiter|grant[8]~q ),
	.asdata(vcc),
	.clrn(resync_chains0sync_r_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reg_grant_last[8]~q ),
	.prn(vcc));
defparam \reg_grant_last[8] .is_wysiwyg = "true";
defparam \reg_grant_last[8] .power_up = "low";

cyclonev_lcell_comb \lif_is_active~0 (
	.dataa(!\arbiter|grant[7]~q ),
	.datab(!\arbiter|grant[8]~q ),
	.datac(!\reg_grant_last[7]~q ),
	.datad(!\reg_grant_last[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_is_active~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_is_active~0 .extended_lut = "off";
defparam \lif_is_active~0 .lut_mask = 64'h8421842184218421;
defparam \lif_is_active~0 .shared_arith = "off";

dffeas \reg_grant_last[0] (
	.clk(mgmt_clk_clk),
	.d(\arbiter|grant[0]~q ),
	.asdata(vcc),
	.clrn(resync_chains0sync_r_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reg_grant_last[0]~q ),
	.prn(vcc));
defparam \reg_grant_last[0] .is_wysiwyg = "true";
defparam \reg_grant_last[0] .power_up = "low";

dffeas \reg_grant_last[1] (
	.clk(mgmt_clk_clk),
	.d(\arbiter|grant[1]~q ),
	.asdata(vcc),
	.clrn(resync_chains0sync_r_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reg_grant_last[1]~q ),
	.prn(vcc));
defparam \reg_grant_last[1] .is_wysiwyg = "true";
defparam \reg_grant_last[1] .power_up = "low";

cyclonev_lcell_comb \lif_is_active~1 (
	.dataa(!\arbiter|grant[0]~q ),
	.datab(!\arbiter|grant[1]~q ),
	.datac(!\reg_grant_last[0]~q ),
	.datad(!\reg_grant_last[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_is_active~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_is_active~1 .extended_lut = "off";
defparam \lif_is_active~1 .lut_mask = 64'h8421842184218421;
defparam \lif_is_active~1 .shared_arith = "off";

cyclonev_lcell_comb lif_is_active(
	.dataa(!\arbiter|grant[4]~q ),
	.datab(!\arbiter|WideNor0~combout ),
	.datac(!\reg_grant_last[4]~q ),
	.datad(!\lif_is_active~0_combout ),
	.datae(!\lif_is_active~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_is_active~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam lif_is_active.extended_lut = "off";
defparam lif_is_active.lut_mask = 64'h0000002100000021;
defparam lif_is_active.shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][0] (
	.dataa(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[0]~q ),
	.datab(!\Equal3~0_combout ),
	.datac(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[0]~q ),
	.datad(!\Equal4~0_combout ),
	.datae(!\wmgmt_readdata[8][0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_0_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][0] .extended_lut = "off";
defparam \wmgmt_readdata[8][0] .lut_mask = 64'h111FFFFF111FFFFF;
defparam \wmgmt_readdata[8][0] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][1] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[1]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[1]~q ),
	.datae(!\wmgmt_readdata[8][1]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_1_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][1] .extended_lut = "off";
defparam \wmgmt_readdata[8][1] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][1] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][2] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[2]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[2]~q ),
	.datae(!\wmgmt_readdata[8][2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_2_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][2] .extended_lut = "off";
defparam \wmgmt_readdata[8][2] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][2] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][3] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[3]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[3]~q ),
	.datae(!\wmgmt_readdata[8][3]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_3_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][3] .extended_lut = "off";
defparam \wmgmt_readdata[8][3] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][3] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][4] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[4]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[4]~q ),
	.datae(!\wmgmt_readdata[8][4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_4_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][4] .extended_lut = "off";
defparam \wmgmt_readdata[8][4] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][4] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][5] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[5]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[5]~q ),
	.datae(!\wmgmt_readdata[8][5]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_5_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][5] .extended_lut = "off";
defparam \wmgmt_readdata[8][5] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][5] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][6] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[6]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[6]~q ),
	.datae(!\wmgmt_readdata[8][6]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_6_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][6] .extended_lut = "off";
defparam \wmgmt_readdata[8][6] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][6] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][7] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[7]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[7]~q ),
	.datae(!\wmgmt_readdata[8][7]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_7_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][7] .extended_lut = "off";
defparam \wmgmt_readdata[8][7] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][7] .shared_arith = "off";

cyclonev_lcell_comb \reconfig_mgmt_readdata[8]~3 (
	.dataa(!reconfig_busy),
	.datab(!\Equal4~0_combout ),
	.datac(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[8]~q ),
	.datad(!\reconfig_mgmt_readdata[8]~0_combout ),
	.datae(!\reconfig_mgmt_readdata[8]~1_combout ),
	.dataf(!\reconfig_mgmt_readdata[8]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reconfig_mgmt_readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \reconfig_mgmt_readdata[8]~3 .extended_lut = "off";
defparam \reconfig_mgmt_readdata[8]~3 .lut_mask = 64'h03ABFFFFFFFFFFFF;
defparam \reconfig_mgmt_readdata[8]~3 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][9] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[9]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[9]~q ),
	.datae(!\wmgmt_readdata[8][9]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_9_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][9] .extended_lut = "off";
defparam \wmgmt_readdata[8][9] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][9] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][10] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[10]~q ),
	.datad(!\wmgmt_readdata~9_combout ),
	.datae(!\wmgmt_readdata~10_combout ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_10_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][10] .extended_lut = "off";
defparam \wmgmt_readdata[8][10] .lut_mask = 64'h05FFFFFF37FFFFFF;
defparam \wmgmt_readdata[8][10] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][11] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[11]~q ),
	.datad(!\wmgmt_readdata~11_combout ),
	.datae(!\wmgmt_readdata~12_combout ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_11_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][11] .extended_lut = "off";
defparam \wmgmt_readdata[8][11] .lut_mask = 64'h05FFFFFF37FFFFFF;
defparam \wmgmt_readdata[8][11] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][12] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[12]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[12]~q ),
	.datae(!\wmgmt_readdata[8][12]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_12_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][12] .extended_lut = "off";
defparam \wmgmt_readdata[8][12] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][12] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][13] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[13]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[13]~q ),
	.datae(!\wmgmt_readdata[8][13]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_13_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][13] .extended_lut = "off";
defparam \wmgmt_readdata[8][13] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][13] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][14] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[14]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[14]~q ),
	.datae(!\wmgmt_readdata[8][14]~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_14_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][14] .extended_lut = "off";
defparam \wmgmt_readdata[8][14] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][14] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][15] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[15]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[15]~q ),
	.datae(!\wmgmt_readdata[8][15]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_15_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][15] .extended_lut = "off";
defparam \wmgmt_readdata[8][15] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][15] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][16] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[16]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[16]~q ),
	.datae(!\wmgmt_readdata[8][16]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_16_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][16] .extended_lut = "off";
defparam \wmgmt_readdata[8][16] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][16] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][17] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[17]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[17]~q ),
	.datae(!\wmgmt_readdata[8][17]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_17_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][17] .extended_lut = "off";
defparam \wmgmt_readdata[8][17] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][17] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][18] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[18]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[18]~q ),
	.datae(!\wmgmt_readdata[8][18]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_18_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][18] .extended_lut = "off";
defparam \wmgmt_readdata[8][18] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][18] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][19] (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[19]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[19]~q ),
	.datae(!\wmgmt_readdata[8][19]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_19_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][19] .extended_lut = "off";
defparam \wmgmt_readdata[8][19] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][19] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][20] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[20]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[20]~q ),
	.datae(!\wmgmt_readdata[8][20]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_20_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][20] .extended_lut = "off";
defparam \wmgmt_readdata[8][20] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][20] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][21] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[21]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[21]~q ),
	.datae(!\wmgmt_readdata[8][21]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_21_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][21] .extended_lut = "off";
defparam \wmgmt_readdata[8][21] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][21] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][22] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[22]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[22]~q ),
	.datae(!\wmgmt_readdata[8][22]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_22_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][22] .extended_lut = "off";
defparam \wmgmt_readdata[8][22] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][22] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][23] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[23]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[23]~q ),
	.datae(!\wmgmt_readdata[8][23]~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_23_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][23] .extended_lut = "off";
defparam \wmgmt_readdata[8][23] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][23] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][24] (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[24]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[24]~q ),
	.datae(!\wmgmt_readdata[8][24]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_24_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][24] .extended_lut = "off";
defparam \wmgmt_readdata[8][24] .lut_mask = 64'h0537FFFF0537FFFF;
defparam \wmgmt_readdata[8][24] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][25] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(!\wmgmt_readdata~26_combout ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[25]~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[25]~q ),
	.dataf(!\wmgmt_readdata~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_25_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][25] .extended_lut = "off";
defparam \wmgmt_readdata[8][25] .lut_mask = 64'h0F5F3F7FFFFFFFFF;
defparam \wmgmt_readdata[8][25] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][26] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(!\wmgmt_readdata~28_combout ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[26]~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[26]~q ),
	.dataf(!\wmgmt_readdata~29_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_26_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][26] .extended_lut = "off";
defparam \wmgmt_readdata[8][26] .lut_mask = 64'h0F5F3F7FFFFFFFFF;
defparam \wmgmt_readdata[8][26] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][27] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(!\wmgmt_readdata~30_combout ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[27]~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[27]~q ),
	.dataf(!\wmgmt_readdata~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_27_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][27] .extended_lut = "off";
defparam \wmgmt_readdata[8][27] .lut_mask = 64'h0F5F3F7FFFFFFFFF;
defparam \wmgmt_readdata[8][27] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][28] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(!\wmgmt_readdata~32_combout ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[28]~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[28]~q ),
	.dataf(!\wmgmt_readdata~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_28_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][28] .extended_lut = "off";
defparam \wmgmt_readdata[8][28] .lut_mask = 64'h0F5F3F7FFFFFFFFF;
defparam \wmgmt_readdata[8][28] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][29] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(!\wmgmt_readdata~34_combout ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[29]~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[29]~q ),
	.dataf(!\wmgmt_readdata~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_29_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][29] .extended_lut = "off";
defparam \wmgmt_readdata[8][29] .lut_mask = 64'h0F5F3F7FFFFFFFFF;
defparam \wmgmt_readdata[8][29] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][30] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(!\wmgmt_readdata~36_combout ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[30]~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[30]~q ),
	.dataf(!\wmgmt_readdata~37_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_30_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][30] .extended_lut = "off";
defparam \wmgmt_readdata[8][30] .lut_mask = 64'h0F5F3F7FFFFFFFFF;
defparam \wmgmt_readdata[8][30] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][31] (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(!\wmgmt_readdata~38_combout ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[31]~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[31]~q ),
	.dataf(!\wmgmt_readdata~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_readdata_31_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][31] .extended_lut = "off";
defparam \wmgmt_readdata[8][31] .lut_mask = 64'h0F5F3F7FFFFFFFFF;
defparam \wmgmt_readdata[8][31] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_waitrequest[8]~3 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\direct.sc_direct|reg_arb_req~q ),
	.datac(!\arbiter|grant[4]~q ),
	.datad(!\basic|a5|lif[0].logical_if|lif_csr|lif_waitrequest~1_combout ),
	.datae(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_waitrequest~1_combout ),
	.dataf(!\wmgmt_waitrequest[8]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wmgmt_waitrequest_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_waitrequest[8]~3 .extended_lut = "off";
defparam \wmgmt_waitrequest[8]~3 .lut_mask = 64'hFFFFFFFF11111011;
defparam \wmgmt_waitrequest[8]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h0100010001000100;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h0080008000800080;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][0]~0 (
	.dataa(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[0]~q ),
	.datab(!reconfig_mgmt_address_3),
	.datac(!reconfig_mgmt_address_4),
	.datad(!reconfig_mgmt_address_5),
	.datae(!reconfig_mgmt_address_6),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][0]~0 .extended_lut = "off";
defparam \wmgmt_readdata[8][0]~0 .lut_mask = 64'h1000000010C00000;
defparam \wmgmt_readdata[8][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][1]~1 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[1]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][1]~1 .extended_lut = "off";
defparam \wmgmt_readdata[8][1]~1 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][1]~1 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][2]~2 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[2]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][2]~2 .extended_lut = "off";
defparam \wmgmt_readdata[8][2]~2 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][2]~2 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][3]~3 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[3]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][3]~3 .extended_lut = "off";
defparam \wmgmt_readdata[8][3]~3 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][3]~3 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][4]~4 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[4]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][4]~4 .extended_lut = "off";
defparam \wmgmt_readdata[8][4]~4 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][4]~4 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][5]~5 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[5]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][5]~5 .extended_lut = "off";
defparam \wmgmt_readdata[8][5]~5 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][5]~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h4000400040004000;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h0800080008000800;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][6]~6 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[6]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][6]~6 .extended_lut = "off";
defparam \wmgmt_readdata[8][6]~6 .lut_mask = 64'h0000010000800180;
defparam \wmgmt_readdata[8][6]~6 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][7]~7 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[7]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][7]~7 .extended_lut = "off";
defparam \wmgmt_readdata[8][7]~7 .lut_mask = 64'h0000010000800180;
defparam \wmgmt_readdata[8][7]~7 .shared_arith = "off";

cyclonev_lcell_comb \reconfig_mgmt_readdata[8]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reconfig_mgmt_readdata[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reconfig_mgmt_readdata[8]~0 .extended_lut = "off";
defparam \reconfig_mgmt_readdata[8]~0 .lut_mask = 64'h4040404040404040;
defparam \reconfig_mgmt_readdata[8]~0 .shared_arith = "off";

cyclonev_lcell_comb \reconfig_mgmt_readdata[8]~1 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\offset.sc_offset|offset_cancellation_av|offset_cancellation_readdata[8]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reconfig_mgmt_readdata[8]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reconfig_mgmt_readdata[8]~1 .extended_lut = "off";
defparam \reconfig_mgmt_readdata[8]~1 .lut_mask = 64'h0000800008008800;
defparam \reconfig_mgmt_readdata[8]~1 .shared_arith = "off";

cyclonev_lcell_comb \reconfig_mgmt_readdata[8]~2 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[8]~q ),
	.dataf(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reconfig_mgmt_readdata[8]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reconfig_mgmt_readdata[8]~2 .extended_lut = "off";
defparam \reconfig_mgmt_readdata[8]~2 .lut_mask = 64'h0000400001004100;
defparam \reconfig_mgmt_readdata[8]~2 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][9]~8 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[9]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][9]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][9]~8 .extended_lut = "off";
defparam \wmgmt_readdata[8][9]~8 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][9]~8 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~9 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~9 .extended_lut = "off";
defparam \wmgmt_readdata~9 .lut_mask = 64'h0000080000000800;
defparam \wmgmt_readdata~9 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~10 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~10 .extended_lut = "off";
defparam \wmgmt_readdata~10 .lut_mask = 64'h0000010000000100;
defparam \wmgmt_readdata~10 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~11 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~11 .extended_lut = "off";
defparam \wmgmt_readdata~11 .lut_mask = 64'h0000080000000800;
defparam \wmgmt_readdata~11 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~12 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~12 .extended_lut = "off";
defparam \wmgmt_readdata~12 .lut_mask = 64'h0000010000000100;
defparam \wmgmt_readdata~12 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][12]~13 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[12]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][12]~13 .extended_lut = "off";
defparam \wmgmt_readdata[8][12]~13 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][12]~13 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][13]~14 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[13]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[13]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][13]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][13]~14 .extended_lut = "off";
defparam \wmgmt_readdata[8][13]~14 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][13]~14 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][14]~15 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[14]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][14]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][14]~15 .extended_lut = "off";
defparam \wmgmt_readdata[8][14]~15 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][14]~15 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][15]~16 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[15]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][15]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][15]~16 .extended_lut = "off";
defparam \wmgmt_readdata[8][15]~16 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][15]~16 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][16]~17 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[16]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][16]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][16]~17 .extended_lut = "off";
defparam \wmgmt_readdata[8][16]~17 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][16]~17 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][17]~18 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[17]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][17]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][17]~18 .extended_lut = "off";
defparam \wmgmt_readdata[8][17]~18 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][17]~18 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][18]~19 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[18]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][18]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][18]~19 .extended_lut = "off";
defparam \wmgmt_readdata[8][18]~19 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][18]~19 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][19]~20 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[19]~q ),
	.dataf(!\basic|a5|lif[0].logical_if|lif_csr|basic_reconfig_readdata[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][19]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][19]~20 .extended_lut = "off";
defparam \wmgmt_readdata[8][19]~20 .lut_mask = 64'h0000400008004800;
defparam \wmgmt_readdata[8][19]~20 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][20]~21 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[20]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][20]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][20]~21 .extended_lut = "off";
defparam \wmgmt_readdata[8][20]~21 .lut_mask = 64'h0000010000800180;
defparam \wmgmt_readdata[8][20]~21 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][21]~22 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[21]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][21]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][21]~22 .extended_lut = "off";
defparam \wmgmt_readdata[8][21]~22 .lut_mask = 64'h0000010000800180;
defparam \wmgmt_readdata[8][21]~22 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][22]~23 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[22]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][22]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][22]~23 .extended_lut = "off";
defparam \wmgmt_readdata[8][22]~23 .lut_mask = 64'h0000010000800180;
defparam \wmgmt_readdata[8][22]~23 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][23]~24 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[23]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][23]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][23]~24 .extended_lut = "off";
defparam \wmgmt_readdata[8][23]~24 .lut_mask = 64'h0000010000800180;
defparam \wmgmt_readdata[8][23]~24 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata[8][24]~25 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|user_reconfig_readdata[24]~q ),
	.dataf(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata[8][24]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata[8][24]~25 .extended_lut = "off";
defparam \wmgmt_readdata[8][24]~25 .lut_mask = 64'h0000010000800180;
defparam \wmgmt_readdata[8][24]~25 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~26 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~26 .extended_lut = "off";
defparam \wmgmt_readdata~26 .lut_mask = 64'h0000400000004000;
defparam \wmgmt_readdata~26 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~27 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~27 .extended_lut = "off";
defparam \wmgmt_readdata~27 .lut_mask = 64'h0000008000000080;
defparam \wmgmt_readdata~27 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~28 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~28 .extended_lut = "off";
defparam \wmgmt_readdata~28 .lut_mask = 64'h0000400000004000;
defparam \wmgmt_readdata~28 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~29 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~29 .extended_lut = "off";
defparam \wmgmt_readdata~29 .lut_mask = 64'h0000008000000080;
defparam \wmgmt_readdata~29 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~30 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~30 .extended_lut = "off";
defparam \wmgmt_readdata~30 .lut_mask = 64'h0000400000004000;
defparam \wmgmt_readdata~30 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~31 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~31 .extended_lut = "off";
defparam \wmgmt_readdata~31 .lut_mask = 64'h0000008000000080;
defparam \wmgmt_readdata~31 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~32 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~32 .extended_lut = "off";
defparam \wmgmt_readdata~32 .lut_mask = 64'h0000400000004000;
defparam \wmgmt_readdata~32 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~33 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~33 .extended_lut = "off";
defparam \wmgmt_readdata~33 .lut_mask = 64'h0000008000000080;
defparam \wmgmt_readdata~33 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~34 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~34 .extended_lut = "off";
defparam \wmgmt_readdata~34 .lut_mask = 64'h0000400000004000;
defparam \wmgmt_readdata~34 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~35 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~35 .extended_lut = "off";
defparam \wmgmt_readdata~35 .lut_mask = 64'h0000008000000080;
defparam \wmgmt_readdata~35 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~36 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~36 .extended_lut = "off";
defparam \wmgmt_readdata~36 .lut_mask = 64'h0000400000004000;
defparam \wmgmt_readdata~36 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~37 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~37 .extended_lut = "off";
defparam \wmgmt_readdata~37 .lut_mask = 64'h0000008000000080;
defparam \wmgmt_readdata~37 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~38 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|user_reconfig_readdata[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~38 .extended_lut = "off";
defparam \wmgmt_readdata~38 .lut_mask = 64'h0000400000004000;
defparam \wmgmt_readdata~38 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_readdata~39 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|user_reconfig_readdata[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_readdata~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_readdata~39 .extended_lut = "off";
defparam \wmgmt_readdata~39 .lut_mask = 64'h0000008000000080;
defparam \wmgmt_readdata~39 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h8000800080008000;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_waitrequest[0] (
	.dataa(!\Equal0~0_combout ),
	.datab(!\offset.sc_offset|offset_cancellation_av|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ),
	.datac(!reconfig_mgmt_read),
	.datad(!\offset.sc_offset|offset_cancellation_av|wait_gen|launch_reg~q ),
	.datae(!\offset.sc_offset|offset_cancellation_av|wait_gen|wait_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_waitrequest[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_waitrequest[0] .extended_lut = "off";
defparam \wmgmt_waitrequest[0] .lut_mask = 64'h4544454545444545;
defparam \wmgmt_waitrequest[0] .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_waitrequest~0 (
	.dataa(!\Equal3~0_combout ),
	.datab(!reconfig_mgmt_read),
	.datac(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ),
	.datad(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|launch_reg~q ),
	.datae(!\mif.sc_mif|mif_strm_av|inst_xreconf_uif|wait_gen|wait_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_waitrequest~0 .extended_lut = "off";
defparam \wmgmt_waitrequest~0 .lut_mask = 64'h5150515151505151;
defparam \wmgmt_waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_waitrequest~1 (
	.dataa(!\Equal4~0_combout ),
	.datab(!reconfig_mgmt_read),
	.datac(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|rst_sync|resync_chains[0].sync_r[1]~q ),
	.datad(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|launch_reg~q ),
	.datae(!\pll.sc_pll|pll_reconfig_av|inst_pll_uif|wait_gen|wait_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_waitrequest~1 .extended_lut = "off";
defparam \wmgmt_waitrequest~1 .lut_mask = 64'h5150515151505151;
defparam \wmgmt_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \wmgmt_waitrequest[8]~2 (
	.dataa(!\Equal1~0_combout ),
	.datab(!\wmgmt_waitrequest[0]~combout ),
	.datac(!\analog.sc_analog|reconfig_analog_cv|inst_xreconf_uif|wait_gen|wait_req~0_combout ),
	.datad(!\wmgmt_waitrequest~0_combout ),
	.datae(!\wmgmt_waitrequest~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wmgmt_waitrequest[8]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wmgmt_waitrequest[8]~2 .extended_lut = "off";
defparam \wmgmt_waitrequest[8]~2 .lut_mask = 64'h8C0000008C000000;
defparam \wmgmt_waitrequest[8]~2 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_arbiter (
	reg_arb_req,
	grant_4,
	mutex_grant,
	grant_0,
	req_and_use_mutex,
	grant_1,
	mutex_req,
	grant_7,
	mutex_req1,
	grant_8,
	mutex_req2,
	mutex_grant1,
	mutex_grant2,
	mutex_grant3,
	WideNor01,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	reg_arb_req;
output 	grant_4;
input 	mutex_grant;
output 	grant_0;
input 	req_and_use_mutex;
output 	grant_1;
input 	mutex_req;
output 	grant_7;
input 	mutex_req1;
output 	grant_8;
input 	mutex_req2;
input 	mutex_grant1;
input 	mutex_grant2;
input 	mutex_grant3;
output 	WideNor01;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \grant~0_combout ;
wire \grant~2_combout ;
wire \grant~6_combout ;
wire \grant~3_combout ;
wire \grant~1_combout ;
wire \grant~4_combout ;
wire \grant~5_combout ;


dffeas \grant[4] (
	.clk(mgmt_clk_clk),
	.d(\grant~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(grant_4),
	.prn(vcc));
defparam \grant[4] .is_wysiwyg = "true";
defparam \grant[4] .power_up = "low";

dffeas \grant[0] (
	.clk(mgmt_clk_clk),
	.d(\grant~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(grant_0),
	.prn(vcc));
defparam \grant[0] .is_wysiwyg = "true";
defparam \grant[0] .power_up = "low";

dffeas \grant[1] (
	.clk(mgmt_clk_clk),
	.d(\grant~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(grant_1),
	.prn(vcc));
defparam \grant[1] .is_wysiwyg = "true";
defparam \grant[1] .power_up = "low";

dffeas \grant[7] (
	.clk(mgmt_clk_clk),
	.d(\grant~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(grant_7),
	.prn(vcc));
defparam \grant[7] .is_wysiwyg = "true";
defparam \grant[7] .power_up = "low";

dffeas \grant[8] (
	.clk(mgmt_clk_clk),
	.d(\grant~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(grant_8),
	.prn(vcc));
defparam \grant[8] .is_wysiwyg = "true";
defparam \grant[8] .power_up = "low";

cyclonev_lcell_comb WideNor0(
	.dataa(!mutex_req1),
	.datab(!mutex_req2),
	.datac(!\grant~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideNor01),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor0.extended_lut = "off";
defparam WideNor0.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam WideNor0.shared_arith = "off";

cyclonev_lcell_comb \grant~0 (
	.dataa(!req_and_use_mutex),
	.datab(!mutex_grant1),
	.datac(!mutex_grant3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant~0 .extended_lut = "off";
defparam \grant~0 .lut_mask = 64'h8080808080808080;
defparam \grant~0 .shared_arith = "off";

cyclonev_lcell_comb \grant~2 (
	.dataa(!reg_arb_req),
	.datab(!grant_4),
	.datac(!mutex_req),
	.datad(!\grant~0_combout ),
	.datae(!WideNor01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant~2 .extended_lut = "off";
defparam \grant~2 .lut_mask = 64'h3373115133731151;
defparam \grant~2 .shared_arith = "off";

cyclonev_lcell_comb \grant~6 (
	.dataa(!mutex_grant3),
	.datab(!mutex_grant1),
	.datac(!mutex_grant),
	.datad(!mutex_grant2),
	.datae(!req_and_use_mutex),
	.dataf(!grant_0),
	.datag(!WideNor01),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant~6 .extended_lut = "on";
defparam \grant~6 .lut_mask = 64'h00008000F0F0FFFF;
defparam \grant~6 .shared_arith = "off";

cyclonev_lcell_comb \grant~3 (
	.dataa(!mutex_grant),
	.datab(!grant_1),
	.datac(!mutex_req),
	.datad(!\grant~0_combout ),
	.datae(!WideNor01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant~3 .extended_lut = "off";
defparam \grant~3 .lut_mask = 64'h333B030B333B030B;
defparam \grant~3 .shared_arith = "off";

cyclonev_lcell_comb \grant~1 (
	.dataa(!reg_arb_req),
	.datab(!req_and_use_mutex),
	.datac(!mutex_req),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant~1 .extended_lut = "off";
defparam \grant~1 .lut_mask = 64'h8080808080808080;
defparam \grant~1 .shared_arith = "off";

cyclonev_lcell_comb \grant~4 (
	.dataa(!grant_7),
	.datab(!mutex_req1),
	.datac(!grant_8),
	.datad(!mutex_req2),
	.datae(!\grant~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant~4 .extended_lut = "off";
defparam \grant~4 .lut_mask = 64'h1111773111117731;
defparam \grant~4 .shared_arith = "off";

cyclonev_lcell_comb \grant~5 (
	.dataa(!mutex_req1),
	.datab(!grant_8),
	.datac(!mutex_req2),
	.datad(!\grant~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant~5 .extended_lut = "off";
defparam \grant~5 .lut_mask = 64'h032B032B032B032B;
defparam \grant~5 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_analog (
	user_reconfig_readdata_6,
	user_reconfig_readdata_7,
	user_reconfig_readdata_10,
	user_reconfig_readdata_11,
	user_reconfig_readdata_12,
	basic_reconfig_readdata_12,
	user_reconfig_readdata_13,
	basic_reconfig_readdata_13,
	user_reconfig_readdata_14,
	basic_reconfig_readdata_14,
	user_reconfig_readdata_15,
	basic_reconfig_readdata_15,
	user_reconfig_readdata_16,
	basic_reconfig_readdata_16,
	user_reconfig_readdata_17,
	basic_reconfig_readdata_17,
	user_reconfig_readdata_18,
	basic_reconfig_readdata_18,
	user_reconfig_readdata_19,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_11,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	rtl,
	user_reconfig_readdata_0,
	basic_reconfig_readdata_0,
	user_reconfig_readdata_1,
	basic_reconfig_readdata_1,
	user_reconfig_readdata_2,
	basic_reconfig_readdata_2,
	user_reconfig_readdata_3,
	basic_reconfig_readdata_3,
	user_reconfig_readdata_4,
	basic_reconfig_readdata_4,
	user_reconfig_readdata_5,
	basic_reconfig_readdata_5,
	Equal1,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	user_reconfig_readdata_8,
	user_reconfig_readdata_9,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	user_reconfig_readdata_20,
	user_reconfig_readdata_21,
	user_reconfig_readdata_22,
	user_reconfig_readdata_23,
	user_reconfig_readdata_24,
	user_reconfig_readdata_25,
	user_reconfig_readdata_26,
	user_reconfig_readdata_27,
	user_reconfig_readdata_28,
	user_reconfig_readdata_29,
	user_reconfig_readdata_30,
	user_reconfig_readdata_31,
	master_write,
	grant_1,
	mutex_req,
	master_address_2,
	mutex_grant,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	comb,
	analog_reconfig_waitrequest,
	stateSTATE_IDLE,
	ifsel_notdone_resync,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_0,
	Decoder3,
	readdata_for_user_2,
	readdata_for_user_0,
	readdata_for_user_3,
	readdata_for_user_1,
	Decoder31,
	Selector2,
	Selector21,
	Decoder32,
	lpbk_lock,
	analog_offset_0,
	readdata_for_user_10,
	readdata_for_user_8,
	readdata_for_user_11,
	readdata_for_user_9,
	rtl1,
	readdata_for_user_6,
	readdata_for_user_4,
	readdata_for_user_7,
	readdata_for_user_5,
	readdata_for_user_14,
	readdata_for_user_12,
	readdata_for_user_15,
	readdata_for_user_13,
	rtl2,
	rtl3,
	rtl4,
	rtl5,
	rtl6,
	readdata_for_user_16,
	rtl7,
	rtl8,
	WideOr4,
	WideOr41,
	analog_length,
	analog_length1,
	analog_length2,
	rtl9,
	readdata_for_user_17,
	rtl10,
	rtl11,
	user_reconfig_readdata_101,
	rtl12,
	readdata_for_user_18,
	rtl13,
	rtl14,
	uif_writedata_4,
	readdata_for_user_19,
	rtl15,
	rtl16,
	LessThan4,
	readdata_for_user_20,
	rtl17,
	rtl18,
	readdata_for_user_21,
	rtl19,
	rtl20,
	readdata_for_user_22,
	rtl21,
	rtl22,
	readdata_for_user_23,
	rtl23,
	readdata_for_user_24,
	rtl24,
	readdata_for_user_25,
	rtl25,
	readdata_for_user_26,
	rtl26,
	readdata_for_user_27,
	rtl27,
	readdata_for_user_28,
	rtl28,
	readdata_for_user_29,
	rtl29,
	readdata_for_user_30,
	rtl30,
	readdata_for_user_31,
	rtl31,
	rtl32,
	rtl33,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	uif_mode_0,
	Mux0,
	Mux3,
	WideOr0,
	Selector5,
	result_data_0,
	rtl34,
	rtl35,
	rtl36,
	rtl37,
	rtl38,
	rtl39,
	rtl40,
	rtl41,
	rtl42,
	rtl43,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_6;
output 	user_reconfig_readdata_7;
output 	user_reconfig_readdata_10;
output 	user_reconfig_readdata_11;
output 	user_reconfig_readdata_12;
input 	basic_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
input 	basic_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
input 	basic_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
input 	basic_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
input 	basic_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
input 	basic_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
input 	basic_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	master_writedata_16;
output 	master_writedata_17;
output 	master_writedata_18;
output 	master_writedata_19;
output 	master_writedata_20;
output 	master_writedata_21;
output 	master_writedata_22;
output 	master_writedata_23;
output 	master_writedata_24;
output 	master_writedata_25;
output 	master_writedata_26;
output 	master_writedata_27;
output 	master_writedata_11;
output 	master_writedata_28;
output 	master_writedata_12;
output 	master_writedata_29;
output 	master_writedata_13;
output 	master_writedata_30;
output 	master_writedata_14;
output 	master_writedata_31;
output 	master_writedata_15;
input 	rtl;
output 	user_reconfig_readdata_0;
input 	basic_reconfig_readdata_0;
output 	user_reconfig_readdata_1;
input 	basic_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
input 	basic_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
input 	basic_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
input 	basic_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
input 	basic_reconfig_readdata_5;
input 	Equal1;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
output 	user_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	user_reconfig_readdata_20;
output 	user_reconfig_readdata_21;
output 	user_reconfig_readdata_22;
output 	user_reconfig_readdata_23;
output 	user_reconfig_readdata_24;
output 	user_reconfig_readdata_25;
output 	user_reconfig_readdata_26;
output 	user_reconfig_readdata_27;
output 	user_reconfig_readdata_28;
output 	user_reconfig_readdata_29;
output 	user_reconfig_readdata_30;
output 	user_reconfig_readdata_31;
output 	master_write;
input 	grant_1;
output 	mutex_req;
output 	master_address_2;
output 	mutex_grant;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	comb;
output 	analog_reconfig_waitrequest;
output 	stateSTATE_IDLE;
input 	ifsel_notdone_resync;
output 	uif_addr_offset_5;
output 	uif_addr_offset_4;
output 	uif_addr_offset_0;
output 	Decoder3;
output 	readdata_for_user_2;
output 	readdata_for_user_0;
output 	readdata_for_user_3;
output 	readdata_for_user_1;
output 	Decoder31;
output 	Selector2;
output 	Selector21;
output 	Decoder32;
output 	lpbk_lock;
output 	analog_offset_0;
output 	readdata_for_user_10;
output 	readdata_for_user_8;
output 	readdata_for_user_11;
output 	readdata_for_user_9;
input 	rtl1;
output 	readdata_for_user_6;
output 	readdata_for_user_4;
output 	readdata_for_user_7;
output 	readdata_for_user_5;
output 	readdata_for_user_14;
output 	readdata_for_user_12;
output 	readdata_for_user_15;
output 	readdata_for_user_13;
input 	rtl2;
input 	rtl3;
input 	rtl4;
input 	rtl5;
input 	rtl6;
output 	readdata_for_user_16;
input 	rtl7;
input 	rtl8;
output 	WideOr4;
output 	WideOr41;
output 	analog_length;
output 	analog_length1;
output 	analog_length2;
input 	rtl9;
output 	readdata_for_user_17;
input 	rtl10;
input 	rtl11;
input 	user_reconfig_readdata_101;
input 	rtl12;
output 	readdata_for_user_18;
input 	rtl13;
input 	rtl14;
output 	uif_writedata_4;
output 	readdata_for_user_19;
input 	rtl15;
input 	rtl16;
output 	LessThan4;
output 	readdata_for_user_20;
input 	rtl17;
input 	rtl18;
output 	readdata_for_user_21;
input 	rtl19;
input 	rtl20;
output 	readdata_for_user_22;
input 	rtl21;
input 	rtl22;
output 	readdata_for_user_23;
input 	rtl23;
output 	readdata_for_user_24;
input 	rtl24;
output 	readdata_for_user_25;
input 	rtl25;
output 	readdata_for_user_26;
input 	rtl26;
output 	readdata_for_user_27;
input 	rtl27;
output 	readdata_for_user_28;
input 	rtl28;
output 	readdata_for_user_29;
input 	rtl29;
output 	readdata_for_user_30;
input 	rtl30;
output 	readdata_for_user_31;
input 	rtl31;
input 	rtl32;
input 	rtl33;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	uif_mode_0;
input 	Mux0;
input 	Mux3;
output 	WideOr0;
output 	Selector5;
output 	result_data_0;
input 	rtl34;
input 	rtl35;
input 	rtl36;
input 	rtl37;
input 	rtl38;
input 	rtl39;
input 	rtl40;
input 	rtl41;
input 	rtl42;
input 	rtl43;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



RECONFIGURE_IP_alt_xcvr_reconfig_analog_av reconfig_analog_cv(
	.user_reconfig_readdata_6(user_reconfig_readdata_6),
	.user_reconfig_readdata_7(user_reconfig_readdata_7),
	.user_reconfig_readdata_10(user_reconfig_readdata_10),
	.user_reconfig_readdata_11(user_reconfig_readdata_11),
	.user_reconfig_readdata_12(user_reconfig_readdata_12),
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.user_reconfig_readdata_13(user_reconfig_readdata_13),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.user_reconfig_readdata_14(user_reconfig_readdata_14),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.user_reconfig_readdata_15(user_reconfig_readdata_15),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.user_reconfig_readdata_16(user_reconfig_readdata_16),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.user_reconfig_readdata_17(user_reconfig_readdata_17),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.user_reconfig_readdata_18(user_reconfig_readdata_18),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.user_reconfig_readdata_19(user_reconfig_readdata_19),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.master_writedata_16(master_writedata_16),
	.master_writedata_17(master_writedata_17),
	.master_writedata_18(master_writedata_18),
	.master_writedata_19(master_writedata_19),
	.master_writedata_20(master_writedata_20),
	.master_writedata_21(master_writedata_21),
	.master_writedata_22(master_writedata_22),
	.master_writedata_23(master_writedata_23),
	.master_writedata_24(master_writedata_24),
	.master_writedata_25(master_writedata_25),
	.master_writedata_26(master_writedata_26),
	.master_writedata_27(master_writedata_27),
	.master_writedata_11(master_writedata_11),
	.master_writedata_28(master_writedata_28),
	.master_writedata_12(master_writedata_12),
	.master_writedata_29(master_writedata_29),
	.master_writedata_13(master_writedata_13),
	.master_writedata_30(master_writedata_30),
	.master_writedata_14(master_writedata_14),
	.master_writedata_31(master_writedata_31),
	.master_writedata_15(master_writedata_15),
	.rtl(rtl),
	.user_reconfig_readdata_0(user_reconfig_readdata_0),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.user_reconfig_readdata_1(user_reconfig_readdata_1),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.user_reconfig_readdata_2(user_reconfig_readdata_2),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.user_reconfig_readdata_3(user_reconfig_readdata_3),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.user_reconfig_readdata_4(user_reconfig_readdata_4),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.user_reconfig_readdata_5(user_reconfig_readdata_5),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.Equal1(Equal1),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.user_reconfig_readdata_8(user_reconfig_readdata_8),
	.user_reconfig_readdata_9(user_reconfig_readdata_9),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.user_reconfig_readdata_20(user_reconfig_readdata_20),
	.user_reconfig_readdata_21(user_reconfig_readdata_21),
	.user_reconfig_readdata_22(user_reconfig_readdata_22),
	.user_reconfig_readdata_23(user_reconfig_readdata_23),
	.user_reconfig_readdata_24(user_reconfig_readdata_24),
	.user_reconfig_readdata_25(user_reconfig_readdata_25),
	.user_reconfig_readdata_26(user_reconfig_readdata_26),
	.user_reconfig_readdata_27(user_reconfig_readdata_27),
	.user_reconfig_readdata_28(user_reconfig_readdata_28),
	.user_reconfig_readdata_29(user_reconfig_readdata_29),
	.user_reconfig_readdata_30(user_reconfig_readdata_30),
	.user_reconfig_readdata_31(user_reconfig_readdata_31),
	.master_write(master_write),
	.grant_1(grant_1),
	.mutex_req(mutex_req),
	.master_address_2(master_address_2),
	.mutex_grant(mutex_grant),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.comb(comb),
	.analog_reconfig_waitrequest(analog_reconfig_waitrequest),
	.stateSTATE_IDLE(stateSTATE_IDLE),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.uif_addr_offset_5(uif_addr_offset_5),
	.uif_addr_offset_4(uif_addr_offset_4),
	.uif_addr_offset_0(uif_addr_offset_0),
	.Decoder3(Decoder3),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_1(readdata_for_user_1),
	.Decoder31(Decoder31),
	.Selector2(Selector2),
	.Selector21(Selector21),
	.Decoder32(Decoder32),
	.lpbk_lock(lpbk_lock),
	.analog_offset_0(analog_offset_0),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_9(readdata_for_user_9),
	.rtl1(rtl1),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_13(readdata_for_user_13),
	.rtl2(rtl2),
	.rtl3(rtl3),
	.rtl4(rtl4),
	.rtl5(rtl5),
	.rtl6(rtl6),
	.readdata_for_user_16(readdata_for_user_16),
	.rtl7(rtl7),
	.rtl8(rtl8),
	.WideOr4(WideOr4),
	.WideOr41(WideOr41),
	.analog_length(analog_length),
	.analog_length1(analog_length1),
	.analog_length2(analog_length2),
	.rtl9(rtl9),
	.readdata_for_user_17(readdata_for_user_17),
	.rtl10(rtl10),
	.rtl11(rtl11),
	.user_reconfig_readdata_101(user_reconfig_readdata_101),
	.rtl12(rtl12),
	.readdata_for_user_18(readdata_for_user_18),
	.rtl13(rtl13),
	.rtl14(rtl14),
	.uif_writedata_4(uif_writedata_4),
	.readdata_for_user_19(readdata_for_user_19),
	.rtl15(rtl15),
	.rtl16(rtl16),
	.LessThan4(LessThan4),
	.readdata_for_user_20(readdata_for_user_20),
	.rtl17(rtl17),
	.rtl18(rtl18),
	.readdata_for_user_21(readdata_for_user_21),
	.rtl19(rtl19),
	.rtl20(rtl20),
	.readdata_for_user_22(readdata_for_user_22),
	.rtl21(rtl21),
	.rtl22(rtl22),
	.readdata_for_user_23(readdata_for_user_23),
	.rtl23(rtl23),
	.readdata_for_user_24(readdata_for_user_24),
	.rtl24(rtl24),
	.readdata_for_user_25(readdata_for_user_25),
	.rtl25(rtl25),
	.readdata_for_user_26(readdata_for_user_26),
	.rtl26(rtl26),
	.readdata_for_user_27(readdata_for_user_27),
	.rtl27(rtl27),
	.readdata_for_user_28(readdata_for_user_28),
	.rtl28(rtl28),
	.readdata_for_user_29(readdata_for_user_29),
	.rtl29(rtl29),
	.readdata_for_user_30(readdata_for_user_30),
	.rtl30(rtl30),
	.readdata_for_user_31(readdata_for_user_31),
	.rtl31(rtl31),
	.rtl32(rtl32),
	.rtl33(rtl33),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.uif_mode_0(uif_mode_0),
	.Mux0(Mux0),
	.Mux3(Mux3),
	.WideOr0(WideOr0),
	.Selector5(Selector5),
	.result_data_0(result_data_0),
	.rtl34(rtl34),
	.rtl35(rtl35),
	.rtl36(rtl36),
	.rtl37(rtl37),
	.rtl38(rtl38),
	.rtl39(rtl39),
	.rtl40(rtl40),
	.rtl41(rtl41),
	.rtl42(rtl42),
	.rtl43(rtl43),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15));

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_analog_av (
	user_reconfig_readdata_6,
	user_reconfig_readdata_7,
	user_reconfig_readdata_10,
	user_reconfig_readdata_11,
	user_reconfig_readdata_12,
	basic_reconfig_readdata_12,
	user_reconfig_readdata_13,
	basic_reconfig_readdata_13,
	user_reconfig_readdata_14,
	basic_reconfig_readdata_14,
	user_reconfig_readdata_15,
	basic_reconfig_readdata_15,
	user_reconfig_readdata_16,
	basic_reconfig_readdata_16,
	user_reconfig_readdata_17,
	basic_reconfig_readdata_17,
	user_reconfig_readdata_18,
	basic_reconfig_readdata_18,
	user_reconfig_readdata_19,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_11,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	rtl,
	user_reconfig_readdata_0,
	basic_reconfig_readdata_0,
	user_reconfig_readdata_1,
	basic_reconfig_readdata_1,
	user_reconfig_readdata_2,
	basic_reconfig_readdata_2,
	user_reconfig_readdata_3,
	basic_reconfig_readdata_3,
	user_reconfig_readdata_4,
	basic_reconfig_readdata_4,
	user_reconfig_readdata_5,
	basic_reconfig_readdata_5,
	Equal1,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	user_reconfig_readdata_8,
	user_reconfig_readdata_9,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	user_reconfig_readdata_20,
	user_reconfig_readdata_21,
	user_reconfig_readdata_22,
	user_reconfig_readdata_23,
	user_reconfig_readdata_24,
	user_reconfig_readdata_25,
	user_reconfig_readdata_26,
	user_reconfig_readdata_27,
	user_reconfig_readdata_28,
	user_reconfig_readdata_29,
	user_reconfig_readdata_30,
	user_reconfig_readdata_31,
	master_write,
	grant_1,
	mutex_req,
	master_address_2,
	mutex_grant,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	comb,
	analog_reconfig_waitrequest,
	stateSTATE_IDLE,
	ifsel_notdone_resync,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_0,
	Decoder3,
	readdata_for_user_2,
	readdata_for_user_0,
	readdata_for_user_3,
	readdata_for_user_1,
	Decoder31,
	Selector2,
	Selector21,
	Decoder32,
	lpbk_lock,
	analog_offset_0,
	readdata_for_user_10,
	readdata_for_user_8,
	readdata_for_user_11,
	readdata_for_user_9,
	rtl1,
	readdata_for_user_6,
	readdata_for_user_4,
	readdata_for_user_7,
	readdata_for_user_5,
	readdata_for_user_14,
	readdata_for_user_12,
	readdata_for_user_15,
	readdata_for_user_13,
	rtl2,
	rtl3,
	rtl4,
	rtl5,
	rtl6,
	readdata_for_user_16,
	rtl7,
	rtl8,
	WideOr4,
	WideOr41,
	analog_length,
	analog_length1,
	analog_length2,
	rtl9,
	readdata_for_user_17,
	rtl10,
	rtl11,
	user_reconfig_readdata_101,
	rtl12,
	readdata_for_user_18,
	rtl13,
	rtl14,
	uif_writedata_4,
	readdata_for_user_19,
	rtl15,
	rtl16,
	LessThan4,
	readdata_for_user_20,
	rtl17,
	rtl18,
	readdata_for_user_21,
	rtl19,
	rtl20,
	readdata_for_user_22,
	rtl21,
	rtl22,
	readdata_for_user_23,
	rtl23,
	readdata_for_user_24,
	rtl24,
	readdata_for_user_25,
	rtl25,
	readdata_for_user_26,
	rtl26,
	readdata_for_user_27,
	rtl27,
	readdata_for_user_28,
	rtl28,
	readdata_for_user_29,
	rtl29,
	readdata_for_user_30,
	rtl30,
	readdata_for_user_31,
	rtl31,
	rtl32,
	rtl33,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	uif_mode_0,
	Mux0,
	Mux3,
	WideOr0,
	Selector5,
	result_data_0,
	rtl34,
	rtl35,
	rtl36,
	rtl37,
	rtl38,
	rtl39,
	rtl40,
	rtl41,
	rtl42,
	rtl43,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_6;
output 	user_reconfig_readdata_7;
output 	user_reconfig_readdata_10;
output 	user_reconfig_readdata_11;
output 	user_reconfig_readdata_12;
input 	basic_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
input 	basic_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
input 	basic_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
input 	basic_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
input 	basic_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
input 	basic_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
input 	basic_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	master_writedata_16;
output 	master_writedata_17;
output 	master_writedata_18;
output 	master_writedata_19;
output 	master_writedata_20;
output 	master_writedata_21;
output 	master_writedata_22;
output 	master_writedata_23;
output 	master_writedata_24;
output 	master_writedata_25;
output 	master_writedata_26;
output 	master_writedata_27;
output 	master_writedata_11;
output 	master_writedata_28;
output 	master_writedata_12;
output 	master_writedata_29;
output 	master_writedata_13;
output 	master_writedata_30;
output 	master_writedata_14;
output 	master_writedata_31;
output 	master_writedata_15;
input 	rtl;
output 	user_reconfig_readdata_0;
input 	basic_reconfig_readdata_0;
output 	user_reconfig_readdata_1;
input 	basic_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
input 	basic_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
input 	basic_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
input 	basic_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
input 	basic_reconfig_readdata_5;
input 	Equal1;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
output 	user_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	user_reconfig_readdata_20;
output 	user_reconfig_readdata_21;
output 	user_reconfig_readdata_22;
output 	user_reconfig_readdata_23;
output 	user_reconfig_readdata_24;
output 	user_reconfig_readdata_25;
output 	user_reconfig_readdata_26;
output 	user_reconfig_readdata_27;
output 	user_reconfig_readdata_28;
output 	user_reconfig_readdata_29;
output 	user_reconfig_readdata_30;
output 	user_reconfig_readdata_31;
output 	master_write;
input 	grant_1;
output 	mutex_req;
output 	master_address_2;
output 	mutex_grant;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	comb;
output 	analog_reconfig_waitrequest;
output 	stateSTATE_IDLE;
input 	ifsel_notdone_resync;
output 	uif_addr_offset_5;
output 	uif_addr_offset_4;
output 	uif_addr_offset_0;
output 	Decoder3;
output 	readdata_for_user_2;
output 	readdata_for_user_0;
output 	readdata_for_user_3;
output 	readdata_for_user_1;
output 	Decoder31;
output 	Selector2;
output 	Selector21;
output 	Decoder32;
output 	lpbk_lock;
output 	analog_offset_0;
output 	readdata_for_user_10;
output 	readdata_for_user_8;
output 	readdata_for_user_11;
output 	readdata_for_user_9;
input 	rtl1;
output 	readdata_for_user_6;
output 	readdata_for_user_4;
output 	readdata_for_user_7;
output 	readdata_for_user_5;
output 	readdata_for_user_14;
output 	readdata_for_user_12;
output 	readdata_for_user_15;
output 	readdata_for_user_13;
input 	rtl2;
input 	rtl3;
input 	rtl4;
input 	rtl5;
input 	rtl6;
output 	readdata_for_user_16;
input 	rtl7;
input 	rtl8;
output 	WideOr4;
output 	WideOr41;
output 	analog_length;
output 	analog_length1;
output 	analog_length2;
input 	rtl9;
output 	readdata_for_user_17;
input 	rtl10;
input 	rtl11;
input 	user_reconfig_readdata_101;
input 	rtl12;
output 	readdata_for_user_18;
input 	rtl13;
input 	rtl14;
output 	uif_writedata_4;
output 	readdata_for_user_19;
input 	rtl15;
input 	rtl16;
output 	LessThan4;
output 	readdata_for_user_20;
input 	rtl17;
input 	rtl18;
output 	readdata_for_user_21;
input 	rtl19;
input 	rtl20;
output 	readdata_for_user_22;
input 	rtl21;
input 	rtl22;
output 	readdata_for_user_23;
input 	rtl23;
output 	readdata_for_user_24;
input 	rtl24;
output 	readdata_for_user_25;
input 	rtl25;
output 	readdata_for_user_26;
input 	rtl26;
output 	readdata_for_user_27;
input 	rtl27;
output 	readdata_for_user_28;
input 	rtl28;
output 	readdata_for_user_29;
input 	rtl29;
output 	readdata_for_user_30;
input 	rtl30;
output 	readdata_for_user_31;
input 	rtl31;
input 	rtl32;
input 	rtl33;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	uif_mode_0;
input 	Mux0;
input 	Mux3;
output 	WideOr0;
output 	Selector5;
output 	result_data_0;
input 	rtl34;
input 	rtl35;
input 	rtl36;
input 	rtl37;
input 	rtl38;
input 	rtl39;
input 	rtl40;
input 	rtl41;
input 	rtl42;
input 	rtl43;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \inst_xreconf_uif|uif_addr_offset[1]~q ;
wire \inst_xreconf_uif|uif_addr_offset[3]~q ;
wire \inst_xreconf_uif|uif_addr_offset[2]~q ;
wire \inst_analog_datactrl|Decoder3~1_combout ;
wire \inst_analog_datactrl|Decoder3~4_combout ;
wire \inst_xreconf_uif|uif_mode[1]~q ;
wire \inst_xreconf_uif|uif_mode[0]~q ;
wire \inst_analog_datactrl|Decoder3~5_combout ;
wire \inst_analog_datactrl|lpbk_done~0_combout ;
wire \inst_xreconf_uif|uif_writedata[0]~q ;
wire \inst_analog_datactrl|lpbk_precdr_reg~q ;
wire \inst_analog_datactrl|lpbk_postcdr_reg~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[0]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ;
wire \inst_xreconf_uif|uif_writedata[1]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[1]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ;
wire \inst_xreconf_uif|uif_writedata[2]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[2]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ;
wire \inst_xreconf_uif|uif_writedata[3]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[3]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[4]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ;
wire \inst_xreconf_uif|uif_writedata[5]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[5]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ;
wire \inst_xreconf_uif|uif_writedata[6]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[6]~q ;
wire \inst_xreconf_uif|user_reconfig_readdata[7]~16_combout ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[7]~q ;
wire \inst_analog_datactrl|Equal6~0_combout ;
wire \inst_xreconf_uif|uif_logical_ch_addr[8]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ;
wire \inst_xreconf_uif|uif_logical_ch_addr[9]~q ;
wire \inst_analog_datactrl|uif_illegal_pch_error~q ;
wire \inst_analog_datactrl|uif_illegal_offset_error~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ;
wire \inst_analog_datactrl|ShiftRight0~0_combout ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ;
wire \inst_analog_datactrl|inst_analog_ctrlsm|ctrl_opcode[1]~q ;
wire \inst_analog_datactrl|inst_analog_ctrlsm|ctrl_opcode[0]~q ;
wire \inst_analog_datactrl|inst_analog_ctrlsm|ctrl_go~q ;
wire \inst_analog_datactrl|inst_analog_ctrlsm|ctrl_lock~q ;
wire \inst_xreconf_uif|uif_go~q ;
wire \inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ;
wire \inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[1]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[2]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[0]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[3]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[16]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[17]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[18]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[19]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[20]~q ;
wire \inst_analog_datactrl|WideOr5~0_combout ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[4]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[21]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[5]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[22]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[6]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[23]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[7]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[24]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[8]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[25]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[9]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[26]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[10]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[27]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[11]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[28]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[12]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[29]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[13]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[30]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[14]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[31]~q ;
wire \inst_analog_datactrl|inst_rmw_sm|outdata[15]~q ;


RECONFIGURE_IP_alt_xreconf_analog_datactrl_av inst_analog_datactrl(
	.rtl(rtl),
	.stateSTATE_IDLE(stateSTATE_IDLE),
	.reset(ifsel_notdone_resync),
	.uif_addr_offset_5(uif_addr_offset_5),
	.uif_addr_offset_4(uif_addr_offset_4),
	.uif_addr_offset_0(uif_addr_offset_0),
	.uif_addr_offset_1(\inst_xreconf_uif|uif_addr_offset[1]~q ),
	.uif_addr_offset_3(\inst_xreconf_uif|uif_addr_offset[3]~q ),
	.uif_addr_offset_2(\inst_xreconf_uif|uif_addr_offset[2]~q ),
	.Decoder3(Decoder3),
	.Decoder31(\inst_analog_datactrl|Decoder3~1_combout ),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_1(readdata_for_user_1),
	.Decoder32(Decoder31),
	.Selector2(Selector2),
	.Selector21(Selector21),
	.Decoder33(Decoder32),
	.lpbk_lock1(lpbk_lock),
	.analog_offset_0(analog_offset_0),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_9(readdata_for_user_9),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_13(readdata_for_user_13),
	.rtl1(rtl3),
	.rtl2(rtl4),
	.readdata_for_user_16(readdata_for_user_16),
	.Decoder34(\inst_analog_datactrl|Decoder3~4_combout ),
	.uif_mode_1(\inst_xreconf_uif|uif_mode[1]~q ),
	.uif_mode_0(\inst_xreconf_uif|uif_mode[0]~q ),
	.Decoder35(\inst_analog_datactrl|Decoder3~5_combout ),
	.WideOr4(WideOr4),
	.WideOr41(WideOr41),
	.analog_length(analog_length),
	.analog_length1(analog_length1),
	.analog_length2(analog_length2),
	.lpbk_done1(\inst_analog_datactrl|lpbk_done~0_combout ),
	.uif_writedata_0(\inst_xreconf_uif|uif_writedata[0]~q ),
	.lpbk_precdr_reg1(\inst_analog_datactrl|lpbk_precdr_reg~q ),
	.lpbk_postcdr_reg1(\inst_analog_datactrl|lpbk_postcdr_reg~q ),
	.uif_writedata_1(\inst_xreconf_uif|uif_writedata[1]~q ),
	.uif_writedata_2(\inst_xreconf_uif|uif_writedata[2]~q ),
	.readdata_for_user_17(readdata_for_user_17),
	.uif_writedata_3(\inst_xreconf_uif|uif_writedata[3]~q ),
	.readdata_for_user_18(readdata_for_user_18),
	.readdata_for_user_19(readdata_for_user_19),
	.LessThan4(LessThan4),
	.uif_writedata_5(\inst_xreconf_uif|uif_writedata[5]~q ),
	.readdata_for_user_20(readdata_for_user_20),
	.uif_writedata_6(\inst_xreconf_uif|uif_writedata[6]~q ),
	.readdata_for_user_21(readdata_for_user_21),
	.user_reconfig_readdata_7(\inst_xreconf_uif|user_reconfig_readdata[7]~16_combout ),
	.readdata_for_user_22(readdata_for_user_22),
	.readdata_for_user_23(readdata_for_user_23),
	.Equal6(\inst_analog_datactrl|Equal6~0_combout ),
	.readdata_for_user_24(readdata_for_user_24),
	.uif_illegal_pch_error1(\inst_analog_datactrl|uif_illegal_pch_error~q ),
	.uif_illegal_offset_error1(\inst_analog_datactrl|uif_illegal_offset_error~q ),
	.readdata_for_user_25(readdata_for_user_25),
	.readdata_for_user_26(readdata_for_user_26),
	.readdata_for_user_27(readdata_for_user_27),
	.readdata_for_user_28(readdata_for_user_28),
	.readdata_for_user_29(readdata_for_user_29),
	.readdata_for_user_30(readdata_for_user_30),
	.readdata_for_user_31(readdata_for_user_31),
	.ShiftRight0(\inst_analog_datactrl|ShiftRight0~0_combout ),
	.ctrl_opcode_1(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_opcode[1]~q ),
	.ctrl_opcode_0(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_opcode[0]~q ),
	.ctrl_go(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_go~q ),
	.ctrl_lock(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_lock~q ),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest2),
	.uif_go(\inst_xreconf_uif|uif_go~q ),
	.waitrequest_to_ctrl(\inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ),
	.illegal_phy_ch(\inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ),
	.outdata_1(\inst_analog_datactrl|inst_rmw_sm|outdata[1]~q ),
	.outdata_2(\inst_analog_datactrl|inst_rmw_sm|outdata[2]~q ),
	.outdata_0(\inst_analog_datactrl|inst_rmw_sm|outdata[0]~q ),
	.outdata_3(\inst_analog_datactrl|inst_rmw_sm|outdata[3]~q ),
	.outdata_16(\inst_analog_datactrl|inst_rmw_sm|outdata[16]~q ),
	.outdata_17(\inst_analog_datactrl|inst_rmw_sm|outdata[17]~q ),
	.outdata_18(\inst_analog_datactrl|inst_rmw_sm|outdata[18]~q ),
	.outdata_19(\inst_analog_datactrl|inst_rmw_sm|outdata[19]~q ),
	.outdata_20(\inst_analog_datactrl|inst_rmw_sm|outdata[20]~q ),
	.WideOr5(\inst_analog_datactrl|WideOr5~0_combout ),
	.outdata_4(\inst_analog_datactrl|inst_rmw_sm|outdata[4]~q ),
	.outdata_21(\inst_analog_datactrl|inst_rmw_sm|outdata[21]~q ),
	.outdata_5(\inst_analog_datactrl|inst_rmw_sm|outdata[5]~q ),
	.outdata_22(\inst_analog_datactrl|inst_rmw_sm|outdata[22]~q ),
	.outdata_6(\inst_analog_datactrl|inst_rmw_sm|outdata[6]~q ),
	.outdata_23(\inst_analog_datactrl|inst_rmw_sm|outdata[23]~q ),
	.outdata_7(\inst_analog_datactrl|inst_rmw_sm|outdata[7]~q ),
	.outdata_24(\inst_analog_datactrl|inst_rmw_sm|outdata[24]~q ),
	.outdata_8(\inst_analog_datactrl|inst_rmw_sm|outdata[8]~q ),
	.outdata_25(\inst_analog_datactrl|inst_rmw_sm|outdata[25]~q ),
	.outdata_9(\inst_analog_datactrl|inst_rmw_sm|outdata[9]~q ),
	.outdata_26(\inst_analog_datactrl|inst_rmw_sm|outdata[26]~q ),
	.outdata_10(\inst_analog_datactrl|inst_rmw_sm|outdata[10]~q ),
	.outdata_27(\inst_analog_datactrl|inst_rmw_sm|outdata[27]~q ),
	.outdata_11(\inst_analog_datactrl|inst_rmw_sm|outdata[11]~q ),
	.outdata_28(\inst_analog_datactrl|inst_rmw_sm|outdata[28]~q ),
	.outdata_12(\inst_analog_datactrl|inst_rmw_sm|outdata[12]~q ),
	.outdata_29(\inst_analog_datactrl|inst_rmw_sm|outdata[29]~q ),
	.outdata_13(\inst_analog_datactrl|inst_rmw_sm|outdata[13]~q ),
	.outdata_30(\inst_analog_datactrl|inst_rmw_sm|outdata[30]~q ),
	.outdata_14(\inst_analog_datactrl|inst_rmw_sm|outdata[14]~q ),
	.outdata_31(\inst_analog_datactrl|inst_rmw_sm|outdata[31]~q ),
	.outdata_15(\inst_analog_datactrl|inst_rmw_sm|outdata[15]~q ),
	.Selector5(Selector5),
	.result_data_0(result_data_0),
	.rtl3(rtl34),
	.rtl4(rtl35),
	.rtl5(rtl36),
	.rtl6(rtl37),
	.rtl7(rtl38),
	.rtl8(rtl39),
	.rtl9(rtl40),
	.rtl10(rtl41),
	.rtl11(rtl42),
	.rtl12(rtl43),
	.clk(mgmt_clk_clk));

RECONFIGURE_IP_alt_xreconf_uif inst_xreconf_uif(
	.user_reconfig_readdata_6(user_reconfig_readdata_6),
	.user_reconfig_readdata_7(user_reconfig_readdata_7),
	.user_reconfig_readdata_10(user_reconfig_readdata_10),
	.user_reconfig_readdata_11(user_reconfig_readdata_11),
	.user_reconfig_readdata_12(user_reconfig_readdata_12),
	.user_reconfig_readdata_13(user_reconfig_readdata_13),
	.user_reconfig_readdata_14(user_reconfig_readdata_14),
	.user_reconfig_readdata_15(user_reconfig_readdata_15),
	.user_reconfig_readdata_16(user_reconfig_readdata_16),
	.user_reconfig_readdata_17(user_reconfig_readdata_17),
	.user_reconfig_readdata_18(user_reconfig_readdata_18),
	.user_reconfig_readdata_19(user_reconfig_readdata_19),
	.user_reconfig_readdata_0(user_reconfig_readdata_0),
	.user_reconfig_readdata_1(user_reconfig_readdata_1),
	.user_reconfig_readdata_2(user_reconfig_readdata_2),
	.user_reconfig_readdata_3(user_reconfig_readdata_3),
	.user_reconfig_readdata_4(user_reconfig_readdata_4),
	.user_reconfig_readdata_5(user_reconfig_readdata_5),
	.Equal1(Equal1),
	.user_reconfig_readdata_8(user_reconfig_readdata_8),
	.user_reconfig_readdata_9(user_reconfig_readdata_9),
	.user_reconfig_readdata_20(user_reconfig_readdata_20),
	.user_reconfig_readdata_21(user_reconfig_readdata_21),
	.user_reconfig_readdata_22(user_reconfig_readdata_22),
	.user_reconfig_readdata_23(user_reconfig_readdata_23),
	.user_reconfig_readdata_24(user_reconfig_readdata_24),
	.user_reconfig_readdata_25(user_reconfig_readdata_25),
	.user_reconfig_readdata_26(user_reconfig_readdata_26),
	.user_reconfig_readdata_27(user_reconfig_readdata_27),
	.user_reconfig_readdata_28(user_reconfig_readdata_28),
	.user_reconfig_readdata_29(user_reconfig_readdata_29),
	.user_reconfig_readdata_30(user_reconfig_readdata_30),
	.user_reconfig_readdata_31(user_reconfig_readdata_31),
	.comb(comb),
	.user_reconfig_waitrequest(analog_reconfig_waitrequest),
	.stateSTATE_IDLE(stateSTATE_IDLE),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.uif_addr_offset_5(uif_addr_offset_5),
	.uif_addr_offset_4(uif_addr_offset_4),
	.uif_addr_offset_0(uif_addr_offset_0),
	.uif_addr_offset_1(\inst_xreconf_uif|uif_addr_offset[1]~q ),
	.uif_addr_offset_3(\inst_xreconf_uif|uif_addr_offset[3]~q ),
	.uif_addr_offset_2(\inst_xreconf_uif|uif_addr_offset[2]~q ),
	.Decoder3(\inst_analog_datactrl|Decoder3~1_combout ),
	.Decoder31(Decoder31),
	.Decoder32(Decoder32),
	.rtl(rtl1),
	.rtl1(rtl2),
	.rtl2(rtl3),
	.rtl3(rtl4),
	.rtl4(rtl5),
	.rtl5(rtl6),
	.rtl6(rtl7),
	.rtl7(rtl8),
	.Decoder33(\inst_analog_datactrl|Decoder3~4_combout ),
	.uif_mode_1(\inst_xreconf_uif|uif_mode[1]~q ),
	.uif_mode_0(\inst_xreconf_uif|uif_mode[0]~q ),
	.Decoder34(\inst_analog_datactrl|Decoder3~5_combout ),
	.WideOr4(WideOr41),
	.analog_length(analog_length),
	.analog_length1(analog_length2),
	.lpbk_done(\inst_analog_datactrl|lpbk_done~0_combout ),
	.uif_writedata_0(\inst_xreconf_uif|uif_writedata[0]~q ),
	.lpbk_precdr_reg(\inst_analog_datactrl|lpbk_precdr_reg~q ),
	.lpbk_postcdr_reg(\inst_analog_datactrl|lpbk_postcdr_reg~q ),
	.uif_logical_ch_addr_0(\inst_xreconf_uif|uif_logical_ch_addr[0]~q ),
	.ph_readdata_0(\inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ),
	.uif_writedata_1(\inst_xreconf_uif|uif_writedata[1]~q ),
	.uif_logical_ch_addr_1(\inst_xreconf_uif|uif_logical_ch_addr[1]~q ),
	.ph_readdata_1(\inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ),
	.uif_writedata_2(\inst_xreconf_uif|uif_writedata[2]~q ),
	.rtl8(rtl9),
	.rtl9(rtl10),
	.rtl10(rtl11),
	.uif_logical_ch_addr_2(\inst_xreconf_uif|uif_logical_ch_addr[2]~q ),
	.ph_readdata_2(\inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ),
	.user_reconfig_readdata_101(user_reconfig_readdata_101),
	.uif_writedata_3(\inst_xreconf_uif|uif_writedata[3]~q ),
	.rtl11(rtl12),
	.rtl12(rtl13),
	.rtl13(rtl14),
	.uif_logical_ch_addr_3(\inst_xreconf_uif|uif_logical_ch_addr[3]~q ),
	.ph_readdata_3(\inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ),
	.uif_writedata_4(uif_writedata_4),
	.rtl14(rtl15),
	.rtl15(rtl16),
	.LessThan4(LessThan4),
	.uif_logical_ch_addr_4(\inst_xreconf_uif|uif_logical_ch_addr[4]~q ),
	.ph_readdata_4(\inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ),
	.uif_writedata_5(\inst_xreconf_uif|uif_writedata[5]~q ),
	.rtl16(rtl17),
	.rtl17(rtl18),
	.uif_logical_ch_addr_5(\inst_xreconf_uif|uif_logical_ch_addr[5]~q ),
	.ph_readdata_5(\inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ),
	.uif_writedata_6(\inst_xreconf_uif|uif_writedata[6]~q ),
	.rtl18(rtl19),
	.rtl19(rtl20),
	.ph_readdata_6(\inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ),
	.uif_logical_ch_addr_6(\inst_xreconf_uif|uif_logical_ch_addr[6]~q ),
	.user_reconfig_readdata_71(\inst_xreconf_uif|user_reconfig_readdata[7]~16_combout ),
	.rtl20(rtl21),
	.rtl21(rtl22),
	.ph_readdata_7(\inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ),
	.uif_logical_ch_addr_7(\inst_xreconf_uif|uif_logical_ch_addr[7]~q ),
	.rtl22(rtl23),
	.Equal6(\inst_analog_datactrl|Equal6~0_combout ),
	.uif_logical_ch_addr_8(\inst_xreconf_uif|uif_logical_ch_addr[8]~q ),
	.ph_readdata_8(\inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ),
	.rtl23(rtl24),
	.ph_readdata_9(\inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ),
	.uif_logical_ch_addr_9(\inst_xreconf_uif|uif_logical_ch_addr[9]~q ),
	.uif_illegal_pch_error(\inst_analog_datactrl|uif_illegal_pch_error~q ),
	.uif_illegal_offset_error(\inst_analog_datactrl|uif_illegal_offset_error~q ),
	.ph_readdata_10(\inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ),
	.rtl24(rtl25),
	.ph_readdata_11(\inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ),
	.rtl25(rtl26),
	.ph_readdata_12(\inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ),
	.rtl26(rtl27),
	.ph_readdata_13(\inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ),
	.rtl27(rtl28),
	.ph_readdata_14(\inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ),
	.rtl28(rtl29),
	.ph_readdata_15(\inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ),
	.rtl29(rtl30),
	.ph_readdata_16(\inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ),
	.rtl30(rtl31),
	.ph_readdata_17(\inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ),
	.rtl31(rtl32),
	.ph_readdata_18(\inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ),
	.rtl32(rtl33),
	.ph_readdata_19(\inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ),
	.ShiftRight0(\inst_analog_datactrl|ShiftRight0~0_combout ),
	.ph_readdata_20(\inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ),
	.ph_readdata_21(\inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ),
	.ph_readdata_22(\inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ),
	.ph_readdata_23(\inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ),
	.ph_readdata_24(\inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ),
	.ph_readdata_25(\inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ),
	.ph_readdata_26(\inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ),
	.ph_readdata_27(\inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ),
	.ph_readdata_28(\inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ),
	.ph_readdata_29(\inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ),
	.ph_readdata_30(\inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ),
	.ph_readdata_31(\inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ),
	.uif_go1(\inst_xreconf_uif|uif_go~q ),
	.uif_mode_01(uif_mode_0),
	.Mux0(Mux0),
	.Mux3(Mux3),
	.WideOr0(WideOr0),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15));

RECONFIGURE_IP_alt_xreconf_cif inst_xreconf_cif(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.master_writedata_16(master_writedata_16),
	.master_writedata_17(master_writedata_17),
	.master_writedata_18(master_writedata_18),
	.master_writedata_19(master_writedata_19),
	.master_writedata_20(master_writedata_20),
	.master_writedata_21(master_writedata_21),
	.master_writedata_22(master_writedata_22),
	.master_writedata_23(master_writedata_23),
	.master_writedata_24(master_writedata_24),
	.master_writedata_25(master_writedata_25),
	.master_writedata_26(master_writedata_26),
	.master_writedata_27(master_writedata_27),
	.master_writedata_11(master_writedata_11),
	.master_writedata_28(master_writedata_28),
	.master_writedata_12(master_writedata_12),
	.master_writedata_29(master_writedata_29),
	.master_writedata_13(master_writedata_13),
	.master_writedata_30(master_writedata_30),
	.master_writedata_14(master_writedata_14),
	.master_writedata_31(master_writedata_31),
	.master_writedata_15(master_writedata_15),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.master_write(master_write),
	.grant_1(grant_1),
	.mutex_req(mutex_req),
	.master_address_2(master_address_2),
	.mutex_grant(mutex_grant),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.uif_addr_offset_5(uif_addr_offset_5),
	.uif_addr_offset_4(uif_addr_offset_4),
	.uif_addr_offset_0(uif_addr_offset_0),
	.uif_addr_offset_1(\inst_xreconf_uif|uif_addr_offset[1]~q ),
	.uif_addr_offset_3(\inst_xreconf_uif|uif_addr_offset[3]~q ),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_1(readdata_for_user_1),
	.Decoder3(Decoder31),
	.lpbk_lock(lpbk_lock),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_9(readdata_for_user_9),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_13(readdata_for_user_13),
	.readdata_for_user_16(readdata_for_user_16),
	.analog_length(analog_length),
	.uif_logical_ch_addr_0(\inst_xreconf_uif|uif_logical_ch_addr[0]~q ),
	.ph_readdata_0(\inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ),
	.uif_logical_ch_addr_1(\inst_xreconf_uif|uif_logical_ch_addr[1]~q ),
	.ph_readdata_1(\inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ),
	.readdata_for_user_17(readdata_for_user_17),
	.uif_logical_ch_addr_2(\inst_xreconf_uif|uif_logical_ch_addr[2]~q ),
	.ph_readdata_2(\inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ),
	.readdata_for_user_18(readdata_for_user_18),
	.uif_logical_ch_addr_3(\inst_xreconf_uif|uif_logical_ch_addr[3]~q ),
	.ph_readdata_3(\inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ),
	.readdata_for_user_19(readdata_for_user_19),
	.uif_logical_ch_addr_4(\inst_xreconf_uif|uif_logical_ch_addr[4]~q ),
	.ph_readdata_4(\inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ),
	.readdata_for_user_20(readdata_for_user_20),
	.uif_logical_ch_addr_5(\inst_xreconf_uif|uif_logical_ch_addr[5]~q ),
	.ph_readdata_5(\inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ),
	.readdata_for_user_21(readdata_for_user_21),
	.ph_readdata_6(\inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ),
	.uif_logical_ch_addr_6(\inst_xreconf_uif|uif_logical_ch_addr[6]~q ),
	.readdata_for_user_22(readdata_for_user_22),
	.ph_readdata_7(\inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ),
	.uif_logical_ch_addr_7(\inst_xreconf_uif|uif_logical_ch_addr[7]~q ),
	.readdata_for_user_23(readdata_for_user_23),
	.uif_logical_ch_addr_8(\inst_xreconf_uif|uif_logical_ch_addr[8]~q ),
	.ph_readdata_8(\inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ),
	.readdata_for_user_24(readdata_for_user_24),
	.ph_readdata_9(\inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ),
	.uif_logical_ch_addr_9(\inst_xreconf_uif|uif_logical_ch_addr[9]~q ),
	.ph_readdata_10(\inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ),
	.readdata_for_user_25(readdata_for_user_25),
	.ph_readdata_11(\inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ),
	.readdata_for_user_26(readdata_for_user_26),
	.ph_readdata_12(\inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ),
	.readdata_for_user_27(readdata_for_user_27),
	.ph_readdata_13(\inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ),
	.readdata_for_user_28(readdata_for_user_28),
	.ph_readdata_14(\inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ),
	.readdata_for_user_29(readdata_for_user_29),
	.ph_readdata_15(\inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ),
	.readdata_for_user_30(readdata_for_user_30),
	.ph_readdata_16(\inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ),
	.readdata_for_user_31(readdata_for_user_31),
	.ph_readdata_17(\inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ),
	.ph_readdata_18(\inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ),
	.ph_readdata_19(\inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ),
	.ph_readdata_20(\inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ),
	.ph_readdata_21(\inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ),
	.ph_readdata_22(\inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ),
	.ph_readdata_23(\inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ),
	.ph_readdata_24(\inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ),
	.ph_readdata_25(\inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ),
	.ph_readdata_26(\inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ),
	.ph_readdata_27(\inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ),
	.ph_readdata_28(\inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ),
	.ph_readdata_29(\inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ),
	.ph_readdata_30(\inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ),
	.ph_readdata_31(\inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.ctrl_opcode_1(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_opcode[1]~q ),
	.ctrl_opcode_0(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_opcode[0]~q ),
	.ctrl_go(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_go~q ),
	.ctrl_lock(\inst_analog_datactrl|inst_analog_ctrlsm|ctrl_lock~q ),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.waitrequest_to_ctrl(\inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ),
	.illegal_phy_ch(\inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ),
	.outdata_1(\inst_analog_datactrl|inst_rmw_sm|outdata[1]~q ),
	.outdata_2(\inst_analog_datactrl|inst_rmw_sm|outdata[2]~q ),
	.outdata_0(\inst_analog_datactrl|inst_rmw_sm|outdata[0]~q ),
	.outdata_3(\inst_analog_datactrl|inst_rmw_sm|outdata[3]~q ),
	.outdata_16(\inst_analog_datactrl|inst_rmw_sm|outdata[16]~q ),
	.outdata_17(\inst_analog_datactrl|inst_rmw_sm|outdata[17]~q ),
	.outdata_18(\inst_analog_datactrl|inst_rmw_sm|outdata[18]~q ),
	.outdata_19(\inst_analog_datactrl|inst_rmw_sm|outdata[19]~q ),
	.outdata_20(\inst_analog_datactrl|inst_rmw_sm|outdata[20]~q ),
	.WideOr5(\inst_analog_datactrl|WideOr5~0_combout ),
	.outdata_4(\inst_analog_datactrl|inst_rmw_sm|outdata[4]~q ),
	.outdata_21(\inst_analog_datactrl|inst_rmw_sm|outdata[21]~q ),
	.outdata_5(\inst_analog_datactrl|inst_rmw_sm|outdata[5]~q ),
	.outdata_22(\inst_analog_datactrl|inst_rmw_sm|outdata[22]~q ),
	.outdata_6(\inst_analog_datactrl|inst_rmw_sm|outdata[6]~q ),
	.outdata_23(\inst_analog_datactrl|inst_rmw_sm|outdata[23]~q ),
	.outdata_7(\inst_analog_datactrl|inst_rmw_sm|outdata[7]~q ),
	.outdata_24(\inst_analog_datactrl|inst_rmw_sm|outdata[24]~q ),
	.outdata_8(\inst_analog_datactrl|inst_rmw_sm|outdata[8]~q ),
	.outdata_25(\inst_analog_datactrl|inst_rmw_sm|outdata[25]~q ),
	.outdata_9(\inst_analog_datactrl|inst_rmw_sm|outdata[9]~q ),
	.outdata_26(\inst_analog_datactrl|inst_rmw_sm|outdata[26]~q ),
	.outdata_10(\inst_analog_datactrl|inst_rmw_sm|outdata[10]~q ),
	.outdata_27(\inst_analog_datactrl|inst_rmw_sm|outdata[27]~q ),
	.outdata_11(\inst_analog_datactrl|inst_rmw_sm|outdata[11]~q ),
	.outdata_28(\inst_analog_datactrl|inst_rmw_sm|outdata[28]~q ),
	.outdata_12(\inst_analog_datactrl|inst_rmw_sm|outdata[12]~q ),
	.outdata_29(\inst_analog_datactrl|inst_rmw_sm|outdata[29]~q ),
	.outdata_13(\inst_analog_datactrl|inst_rmw_sm|outdata[13]~q ),
	.outdata_30(\inst_analog_datactrl|inst_rmw_sm|outdata[30]~q ),
	.outdata_14(\inst_analog_datactrl|inst_rmw_sm|outdata[14]~q ),
	.outdata_31(\inst_analog_datactrl|inst_rmw_sm|outdata[31]~q ),
	.outdata_15(\inst_analog_datactrl|inst_rmw_sm|outdata[15]~q ),
	.mgmt_clk_clk(mgmt_clk_clk));

endmodule

module RECONFIGURE_IP_alt_xreconf_analog_datactrl_av (
	rtl,
	stateSTATE_IDLE,
	reset,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_0,
	uif_addr_offset_1,
	uif_addr_offset_3,
	uif_addr_offset_2,
	Decoder3,
	Decoder31,
	readdata_for_user_2,
	readdata_for_user_0,
	readdata_for_user_3,
	readdata_for_user_1,
	Decoder32,
	Selector2,
	Selector21,
	Decoder33,
	lpbk_lock1,
	analog_offset_0,
	readdata_for_user_10,
	readdata_for_user_8,
	readdata_for_user_11,
	readdata_for_user_9,
	readdata_for_user_6,
	readdata_for_user_4,
	readdata_for_user_7,
	readdata_for_user_5,
	readdata_for_user_14,
	readdata_for_user_12,
	readdata_for_user_15,
	readdata_for_user_13,
	rtl1,
	rtl2,
	readdata_for_user_16,
	Decoder34,
	uif_mode_1,
	uif_mode_0,
	Decoder35,
	WideOr4,
	WideOr41,
	analog_length,
	analog_length1,
	analog_length2,
	lpbk_done1,
	uif_writedata_0,
	lpbk_precdr_reg1,
	lpbk_postcdr_reg1,
	uif_writedata_1,
	uif_writedata_2,
	readdata_for_user_17,
	uif_writedata_3,
	readdata_for_user_18,
	readdata_for_user_19,
	LessThan4,
	uif_writedata_5,
	readdata_for_user_20,
	uif_writedata_6,
	readdata_for_user_21,
	user_reconfig_readdata_7,
	readdata_for_user_22,
	readdata_for_user_23,
	Equal6,
	readdata_for_user_24,
	uif_illegal_pch_error1,
	uif_illegal_offset_error1,
	readdata_for_user_25,
	readdata_for_user_26,
	readdata_for_user_27,
	readdata_for_user_28,
	readdata_for_user_29,
	readdata_for_user_30,
	readdata_for_user_31,
	ShiftRight0,
	ctrl_opcode_1,
	ctrl_opcode_0,
	ctrl_go,
	ctrl_lock,
	basic_reconfig_waitrequest,
	uif_go,
	waitrequest_to_ctrl,
	illegal_phy_ch,
	outdata_1,
	outdata_2,
	outdata_0,
	outdata_3,
	outdata_16,
	outdata_17,
	outdata_18,
	outdata_19,
	outdata_20,
	WideOr5,
	outdata_4,
	outdata_21,
	outdata_5,
	outdata_22,
	outdata_6,
	outdata_23,
	outdata_7,
	outdata_24,
	outdata_8,
	outdata_25,
	outdata_9,
	outdata_26,
	outdata_10,
	outdata_27,
	outdata_11,
	outdata_28,
	outdata_12,
	outdata_29,
	outdata_13,
	outdata_30,
	outdata_14,
	outdata_31,
	outdata_15,
	Selector5,
	result_data_0,
	rtl3,
	rtl4,
	rtl5,
	rtl6,
	rtl7,
	rtl8,
	rtl9,
	rtl10,
	rtl11,
	rtl12,
	clk)/* synthesis synthesis_greybox=0 */;
input 	rtl;
output 	stateSTATE_IDLE;
input 	reset;
input 	uif_addr_offset_5;
input 	uif_addr_offset_4;
input 	uif_addr_offset_0;
input 	uif_addr_offset_1;
input 	uif_addr_offset_3;
input 	uif_addr_offset_2;
output 	Decoder3;
output 	Decoder31;
input 	readdata_for_user_2;
input 	readdata_for_user_0;
input 	readdata_for_user_3;
input 	readdata_for_user_1;
output 	Decoder32;
output 	Selector2;
output 	Selector21;
output 	Decoder33;
output 	lpbk_lock1;
output 	analog_offset_0;
input 	readdata_for_user_10;
input 	readdata_for_user_8;
input 	readdata_for_user_11;
input 	readdata_for_user_9;
input 	readdata_for_user_6;
input 	readdata_for_user_4;
input 	readdata_for_user_7;
input 	readdata_for_user_5;
input 	readdata_for_user_14;
input 	readdata_for_user_12;
input 	readdata_for_user_15;
input 	readdata_for_user_13;
input 	rtl1;
input 	rtl2;
input 	readdata_for_user_16;
output 	Decoder34;
input 	uif_mode_1;
input 	uif_mode_0;
output 	Decoder35;
output 	WideOr4;
output 	WideOr41;
output 	analog_length;
output 	analog_length1;
output 	analog_length2;
output 	lpbk_done1;
input 	uif_writedata_0;
output 	lpbk_precdr_reg1;
output 	lpbk_postcdr_reg1;
input 	uif_writedata_1;
input 	uif_writedata_2;
input 	readdata_for_user_17;
input 	uif_writedata_3;
input 	readdata_for_user_18;
input 	readdata_for_user_19;
output 	LessThan4;
input 	uif_writedata_5;
input 	readdata_for_user_20;
input 	uif_writedata_6;
input 	readdata_for_user_21;
input 	user_reconfig_readdata_7;
input 	readdata_for_user_22;
input 	readdata_for_user_23;
output 	Equal6;
input 	readdata_for_user_24;
output 	uif_illegal_pch_error1;
output 	uif_illegal_offset_error1;
input 	readdata_for_user_25;
input 	readdata_for_user_26;
input 	readdata_for_user_27;
input 	readdata_for_user_28;
input 	readdata_for_user_29;
input 	readdata_for_user_30;
input 	readdata_for_user_31;
output 	ShiftRight0;
output 	ctrl_opcode_1;
output 	ctrl_opcode_0;
output 	ctrl_go;
output 	ctrl_lock;
input 	basic_reconfig_waitrequest;
input 	uif_go;
input 	waitrequest_to_ctrl;
input 	illegal_phy_ch;
output 	outdata_1;
output 	outdata_2;
output 	outdata_0;
output 	outdata_3;
output 	outdata_16;
output 	outdata_17;
output 	outdata_18;
output 	outdata_19;
output 	outdata_20;
output 	WideOr5;
output 	outdata_4;
output 	outdata_21;
output 	outdata_5;
output 	outdata_22;
output 	outdata_6;
output 	outdata_23;
output 	outdata_7;
output 	outdata_24;
output 	outdata_8;
output 	outdata_25;
output 	outdata_9;
output 	outdata_26;
output 	outdata_10;
output 	outdata_27;
output 	outdata_11;
output 	outdata_28;
output 	outdata_12;
output 	outdata_29;
output 	outdata_13;
output 	outdata_30;
output 	outdata_14;
output 	outdata_31;
output 	outdata_15;
output 	Selector5;
output 	result_data_0;
input 	rtl3;
input 	rtl4;
input 	rtl5;
input 	rtl6;
input 	rtl7;
input 	rtl8;
input 	rtl9;
input 	rtl10;
input 	rtl11;
input 	rtl12;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \inst_analog_ctrlsm|lpbk_lock_ack~q ;
wire \lpbk_lock~q ;
wire \lpbk_lock~1_combout ;
wire \Selector6~0_combout ;
wire \Selector6~1_combout ;
wire \lpbk_go~0_combout ;
wire \lpbk_go~q ;
wire \lpbk_done~1_combout ;
wire \lpbk_done~q ;
wire \lpbk_precdr_reg~0_combout ;
wire \lpbk_postcdr_reg~0_combout ;
wire \WideOr11~0_combout ;


RECONFIGURE_IP_alt_xreconf_analog_rmw_av inst_rmw_sm(
	.rtl(rtl),
	.ifsel_notdone_resync(reset),
	.uif_addr_offset_5(uif_addr_offset_5),
	.uif_addr_offset_4(uif_addr_offset_4),
	.uif_addr_offset_1(uif_addr_offset_1),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_1(readdata_for_user_1),
	.Decoder3(Decoder32),
	.Selector2(Selector21),
	.analog_offset_0(analog_offset_0),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_9(readdata_for_user_9),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_13(readdata_for_user_13),
	.rtl1(rtl1),
	.rtl2(rtl2),
	.readdata_for_user_16(readdata_for_user_16),
	.WideOr4(WideOr4),
	.WideOr41(WideOr41),
	.analog_length(analog_length),
	.analog_length1(analog_length1),
	.analog_length2(analog_length2),
	.uif_writedata_2(uif_writedata_2),
	.readdata_for_user_17(readdata_for_user_17),
	.uif_writedata_3(uif_writedata_3),
	.readdata_for_user_18(readdata_for_user_18),
	.readdata_for_user_19(readdata_for_user_19),
	.uif_writedata_5(uif_writedata_5),
	.readdata_for_user_20(readdata_for_user_20),
	.uif_writedata_6(uif_writedata_6),
	.readdata_for_user_21(readdata_for_user_21),
	.readdata_for_user_22(readdata_for_user_22),
	.readdata_for_user_23(readdata_for_user_23),
	.Equal6(Equal6),
	.readdata_for_user_24(readdata_for_user_24),
	.readdata_for_user_25(readdata_for_user_25),
	.readdata_for_user_26(readdata_for_user_26),
	.readdata_for_user_27(readdata_for_user_27),
	.readdata_for_user_28(readdata_for_user_28),
	.readdata_for_user_29(readdata_for_user_29),
	.readdata_for_user_30(readdata_for_user_30),
	.readdata_for_user_31(readdata_for_user_31),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.outdata_1(outdata_1),
	.outdata_2(outdata_2),
	.outdata_0(outdata_0),
	.outdata_3(outdata_3),
	.outdata_16(outdata_16),
	.outdata_17(outdata_17),
	.outdata_18(outdata_18),
	.outdata_19(outdata_19),
	.outdata_20(outdata_20),
	.outdata_4(outdata_4),
	.outdata_21(outdata_21),
	.outdata_5(outdata_5),
	.outdata_22(outdata_22),
	.outdata_6(outdata_6),
	.outdata_23(outdata_23),
	.outdata_7(outdata_7),
	.outdata_24(outdata_24),
	.outdata_8(outdata_8),
	.outdata_25(outdata_25),
	.outdata_9(outdata_9),
	.outdata_26(outdata_26),
	.outdata_10(outdata_10),
	.outdata_27(outdata_27),
	.outdata_11(outdata_11),
	.outdata_28(outdata_28),
	.outdata_12(outdata_12),
	.outdata_29(outdata_29),
	.outdata_13(outdata_13),
	.outdata_30(outdata_30),
	.outdata_14(outdata_14),
	.outdata_31(outdata_31),
	.outdata_15(outdata_15),
	.Selector6(\Selector6~0_combout ),
	.Selector61(\Selector6~1_combout ),
	.result_data_0(result_data_0),
	.rtl3(rtl3),
	.rtl4(rtl4),
	.rtl5(rtl5),
	.rtl6(rtl6),
	.rtl7(rtl7),
	.rtl8(rtl8),
	.rtl9(rtl9),
	.rtl10(rtl10),
	.rtl11(rtl11),
	.rtl12(rtl12),
	.mgmt_clk_clk(clk));

RECONFIGURE_IP_alt_xreconf_analog_ctrlsm inst_analog_ctrlsm(
	.stateSTATE_IDLE(stateSTATE_IDLE),
	.ifsel_notdone_resync(reset),
	.lpbk_lock_ack1(\inst_analog_ctrlsm|lpbk_lock_ack~q ),
	.user_reconfig_readdata_7(user_reconfig_readdata_7),
	.Equal6(Equal6),
	.ctrl_opcode_1(ctrl_opcode_1),
	.ctrl_opcode_0(ctrl_opcode_0),
	.ctrl_go1(ctrl_go),
	.ctrl_lock1(ctrl_lock),
	.uif_go(uif_go),
	.lpbk_go(\lpbk_go~q ),
	.lpbk_lock(\lpbk_lock~q ),
	.waitrequest_to_ctrl(waitrequest_to_ctrl),
	.illegal_phy_ch(illegal_phy_ch),
	.WideOr11(\WideOr11~0_combout ),
	.mgmt_clk_clk(clk));

dffeas lpbk_lock(
	.clk(clk),
	.d(\lpbk_lock~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lpbk_lock~q ),
	.prn(vcc));
defparam lpbk_lock.is_wysiwyg = "true";
defparam lpbk_lock.power_up = "low";

cyclonev_lcell_comb \lpbk_lock~1 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!Decoder3),
	.datae(!lpbk_lock1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpbk_lock~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpbk_lock~1 .extended_lut = "off";
defparam \lpbk_lock~1 .lut_mask = 64'h0000004600000046;
defparam \lpbk_lock~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!uif_addr_offset_0),
	.datab(!lpbk_lock1),
	.datac(!uif_writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \Selector6~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~1 (
	.dataa(!uif_addr_offset_4),
	.datab(!uif_addr_offset_0),
	.datac(!uif_addr_offset_1),
	.datad(!uif_writedata_0),
	.datae(!uif_writedata_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'h00C810D800C810D8;
defparam \Selector6~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder3~0 (
	.dataa(!uif_addr_offset_1),
	.datab(!uif_addr_offset_3),
	.datac(!uif_addr_offset_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder3~0 .extended_lut = "off";
defparam \Decoder3~0 .lut_mask = 64'h8080808080808080;
defparam \Decoder3~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder3~1 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!Decoder3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder3~1 .extended_lut = "off";
defparam \Decoder3~1 .lut_mask = 64'h0004000400040004;
defparam \Decoder3~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder3~2 (
	.dataa(!uif_addr_offset_3),
	.datab(!uif_addr_offset_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder3~2 .extended_lut = "off";
defparam \Decoder3~2 .lut_mask = 64'h8888888888888888;
defparam \Decoder3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!uif_addr_offset_1),
	.datae(!\lpbk_done~q ),
	.dataf(!\inst_analog_ctrlsm|lpbk_lock_ack~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hE680E480E480E480;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!Decoder32),
	.datab(!Selector2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h1111111111111111;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder3~3 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!uif_addr_offset_1),
	.datae(!uif_addr_offset_3),
	.dataf(!uif_addr_offset_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder33),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder3~3 .extended_lut = "off";
defparam \Decoder3~3 .lut_mask = 64'h4000000000000000;
defparam \Decoder3~3 .shared_arith = "off";

cyclonev_lcell_comb \lpbk_lock~0 (
	.dataa(!\lpbk_done~q ),
	.datab(!\inst_analog_ctrlsm|lpbk_lock_ack~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(lpbk_lock1),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpbk_lock~0 .extended_lut = "off";
defparam \lpbk_lock~0 .lut_mask = 64'h8888888888888888;
defparam \lpbk_lock~0 .shared_arith = "off";

cyclonev_lcell_comb \analog_offset[0]~0 (
	.dataa(!Decoder33),
	.datab(!lpbk_lock1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(analog_offset_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \analog_offset[0]~0 .extended_lut = "off";
defparam \analog_offset[0]~0 .lut_mask = 64'h4444444444444444;
defparam \analog_offset[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder3~4 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!Decoder3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder34),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder3~4 .extended_lut = "off";
defparam \Decoder3~4 .lut_mask = 64'h0020002000200020;
defparam \Decoder3~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder3~5 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!uif_addr_offset_1),
	.datae(!Decoder32),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder35),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder3~5 .extended_lut = "off";
defparam \Decoder3~5 .lut_mask = 64'h0000020000000200;
defparam \Decoder3~5 .shared_arith = "off";

cyclonev_lcell_comb \WideOr4~0 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_addr_offset_1),
	.datac(!uif_addr_offset_4),
	.datad(!uif_addr_offset_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr4),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr4~0 .extended_lut = "off";
defparam \WideOr4~0 .lut_mask = 64'h28C028C028C028C0;
defparam \WideOr4~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr4~1 (
	.dataa(!Decoder32),
	.datab(!WideOr4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr41),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr4~1 .extended_lut = "off";
defparam \WideOr4~1 .lut_mask = 64'h1111111111111111;
defparam \WideOr4~1 .shared_arith = "off";

cyclonev_lcell_comb \analog_length~0 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!uif_addr_offset_3),
	.datae(!uif_addr_offset_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(analog_length),
	.sumout(),
	.cout(),
	.shareout());
defparam \analog_length~0 .extended_lut = "off";
defparam \analog_length~0 .lut_mask = 64'h8000000080000000;
defparam \analog_length~0 .shared_arith = "off";

cyclonev_lcell_comb \analog_length~1 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_addr_offset_1),
	.datac(!uif_addr_offset_2),
	.datad(!uif_addr_offset_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(analog_length1),
	.sumout(),
	.cout(),
	.shareout());
defparam \analog_length~1 .extended_lut = "off";
defparam \analog_length~1 .lut_mask = 64'h8040804080408040;
defparam \analog_length~1 .shared_arith = "off";

cyclonev_lcell_comb \analog_length~2 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_3),
	.datac(!analog_length1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(analog_length2),
	.sumout(),
	.cout(),
	.shareout());
defparam \analog_length~2 .extended_lut = "off";
defparam \analog_length~2 .lut_mask = 64'h0808080808080808;
defparam \analog_length~2 .shared_arith = "off";

cyclonev_lcell_comb \lpbk_done~0 (
	.dataa(!Decoder33),
	.datab(!Decoder31),
	.datac(!Decoder35),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(lpbk_done1),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpbk_done~0 .extended_lut = "off";
defparam \lpbk_done~0 .lut_mask = 64'h8080808080808080;
defparam \lpbk_done~0 .shared_arith = "off";

dffeas lpbk_precdr_reg(
	.clk(clk),
	.d(\lpbk_precdr_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lpbk_precdr_reg1),
	.prn(vcc));
defparam lpbk_precdr_reg.is_wysiwyg = "true";
defparam lpbk_precdr_reg.power_up = "low";

dffeas lpbk_postcdr_reg(
	.clk(clk),
	.d(\lpbk_postcdr_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lpbk_postcdr_reg1),
	.prn(vcc));
defparam lpbk_postcdr_reg.is_wysiwyg = "true";
defparam lpbk_postcdr_reg.power_up = "low";

cyclonev_lcell_comb \LessThan4~0 (
	.dataa(!WideOr41),
	.datab(!analog_length),
	.datac(!analog_length2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan4),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~0 .extended_lut = "off";
defparam \LessThan4~0 .lut_mask = 64'h1313131313131313;
defparam \LessThan4~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h2222222222222222;
defparam \Equal6~0 .shared_arith = "off";

dffeas uif_illegal_pch_error(
	.clk(clk),
	.d(illegal_phy_ch),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_illegal_pch_error1),
	.prn(vcc));
defparam uif_illegal_pch_error.is_wysiwyg = "true";
defparam uif_illegal_pch_error.power_up = "low";

dffeas uif_illegal_offset_error(
	.clk(clk),
	.d(\WideOr11~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_illegal_offset_error1),
	.prn(vcc));
defparam uif_illegal_offset_error.is_wysiwyg = "true";
defparam uif_illegal_offset_error.power_up = "low";

cyclonev_lcell_comb \ShiftRight0~0 (
	.dataa(!Decoder32),
	.datab(!Decoder33),
	.datac(!lpbk_lock1),
	.datad(!Selector2),
	.datae(!readdata_for_user_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftRight0),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftRight0~0 .extended_lut = "off";
defparam \ShiftRight0~0 .lut_mask = 64'h0000CF8A0000CF8A;
defparam \ShiftRight0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr5~0 (
	.dataa(!uif_addr_offset_1),
	.datab(!uif_addr_offset_2),
	.datac(!uif_addr_offset_5),
	.datad(!uif_addr_offset_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr5),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr5~0 .extended_lut = "off";
defparam \WideOr5~0 .lut_mask = 64'h0880088008800880;
defparam \WideOr5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!uif_addr_offset_4),
	.datab(!uif_addr_offset_0),
	.datac(!uif_addr_offset_1),
	.datad(!lpbk_lock1),
	.datae(!uif_writedata_0),
	.dataf(!uif_writedata_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h0000001098989898;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \lpbk_go~0 (
	.dataa(!\inst_analog_ctrlsm|lpbk_lock_ack~q ),
	.datab(!lpbk_done1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpbk_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpbk_go~0 .extended_lut = "off";
defparam \lpbk_go~0 .lut_mask = 64'h4444444444444444;
defparam \lpbk_go~0 .shared_arith = "off";

dffeas lpbk_go(
	.clk(clk),
	.d(\lpbk_go~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lpbk_go~q ),
	.prn(vcc));
defparam lpbk_go.is_wysiwyg = "true";
defparam lpbk_go.power_up = "low";

cyclonev_lcell_comb \lpbk_done~1 (
	.dataa(!stateSTATE_IDLE),
	.datab(!\lpbk_done~q ),
	.datac(!\inst_analog_ctrlsm|lpbk_lock_ack~q ),
	.datad(!lpbk_done1),
	.datae(!\lpbk_go~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpbk_done~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpbk_done~1 .extended_lut = "off";
defparam \lpbk_done~1 .lut_mask = 64'h1F003F001F003F00;
defparam \lpbk_done~1 .shared_arith = "off";

dffeas lpbk_done(
	.clk(clk),
	.d(\lpbk_done~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lpbk_done~q ),
	.prn(vcc));
defparam lpbk_done.is_wysiwyg = "true";
defparam lpbk_done.power_up = "low";

cyclonev_lcell_comb \lpbk_precdr_reg~0 (
	.dataa(!lpbk_precdr_reg1),
	.datab(!Decoder33),
	.datac(!Equal6),
	.datad(!uif_writedata_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpbk_precdr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpbk_precdr_reg~0 .extended_lut = "off";
defparam \lpbk_precdr_reg~0 .lut_mask = 64'h5457545754575457;
defparam \lpbk_precdr_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \lpbk_postcdr_reg~0 (
	.dataa(!Equal6),
	.datab(!lpbk_postcdr_reg1),
	.datac(!Decoder31),
	.datad(!uif_writedata_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpbk_postcdr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpbk_postcdr_reg~0 .extended_lut = "off";
defparam \lpbk_postcdr_reg~0 .lut_mask = 64'h3237323732373237;
defparam \lpbk_postcdr_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr11~0 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_1),
	.datad(!uif_addr_offset_0),
	.datae(!uif_addr_offset_2),
	.dataf(!uif_addr_offset_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr11~0 .extended_lut = "off";
defparam \WideOr11~0 .lut_mask = 64'h179FFFFFFFFFFFFF;
defparam \WideOr11~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_analog_ctrlsm (
	stateSTATE_IDLE,
	ifsel_notdone_resync,
	lpbk_lock_ack1,
	user_reconfig_readdata_7,
	Equal6,
	ctrl_opcode_1,
	ctrl_opcode_0,
	ctrl_go1,
	ctrl_lock1,
	uif_go,
	lpbk_go,
	lpbk_lock,
	waitrequest_to_ctrl,
	illegal_phy_ch,
	WideOr11,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	stateSTATE_IDLE;
input 	ifsel_notdone_resync;
output 	lpbk_lock_ack1;
input 	user_reconfig_readdata_7;
input 	Equal6;
output 	ctrl_opcode_1;
output 	ctrl_opcode_0;
output 	ctrl_go1;
output 	ctrl_lock1;
input 	uif_go;
input 	lpbk_go;
input 	lpbk_lock;
input 	waitrequest_to_ctrl;
input 	illegal_phy_ch;
input 	WideOr11;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Selector2~0_combout ;
wire \state.STATE_RMW_GO~q ;
wire \Selector3~0_combout ;
wire \state.STATE_RMW_RD~q ;
wire \next_state.STATE_RMW_WAIT~0_combout ;
wire \state.STATE_RMW_WAIT~q ;
wire \state.STATE_RMW_GO2~q ;
wire \Selector4~0_combout ;
wire \state.STATE_RMW_WR~q ;
wire \next_state.STATE_LOCK_CHK~0_combout ;
wire \state.STATE_LOCK_CHK~q ;
wire \next_state.STATE_GO~0_combout ;
wire \state.STATE_GO~q ;
wire \Selector1~0_combout ;
wire \state.STATE_READ~q ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector5~0_combout ;
wire \ctrl_opcode~0_combout ;
wire \ctrl_opcode~1_combout ;
wire \ctrl_opcode[0]~2_combout ;
wire \ctrl_opcode[0]~3_combout ;
wire \ctrl_go~0_combout ;
wire \ctrl_lock~0_combout ;
wire \ctrl_lock~1_combout ;


dffeas \state.STATE_IDLE (
	.clk(mgmt_clk_clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateSTATE_IDLE),
	.prn(vcc));
defparam \state.STATE_IDLE .is_wysiwyg = "true";
defparam \state.STATE_IDLE .power_up = "low";

dffeas lpbk_lock_ack(
	.clk(mgmt_clk_clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lpbk_lock_ack1),
	.prn(vcc));
defparam lpbk_lock_ack.is_wysiwyg = "true";
defparam lpbk_lock_ack.power_up = "low";

dffeas \ctrl_opcode[1] (
	.clk(mgmt_clk_clk),
	.d(\ctrl_opcode~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_opcode[0]~3_combout ),
	.q(ctrl_opcode_1),
	.prn(vcc));
defparam \ctrl_opcode[1] .is_wysiwyg = "true";
defparam \ctrl_opcode[1] .power_up = "low";

dffeas \ctrl_opcode[0] (
	.clk(mgmt_clk_clk),
	.d(\ctrl_opcode[0]~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_opcode[0]~3_combout ),
	.q(ctrl_opcode_0),
	.prn(vcc));
defparam \ctrl_opcode[0] .is_wysiwyg = "true";
defparam \ctrl_opcode[0] .power_up = "low";

dffeas ctrl_go(
	.clk(mgmt_clk_clk),
	.d(\ctrl_go~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_go1),
	.prn(vcc));
defparam ctrl_go.is_wysiwyg = "true";
defparam ctrl_go.power_up = "low";

dffeas ctrl_lock(
	.clk(mgmt_clk_clk),
	.d(\ctrl_lock~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_lock1),
	.prn(vcc));
defparam ctrl_lock.is_wysiwyg = "true";
defparam ctrl_lock.power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateSTATE_IDLE),
	.datab(!Equal6),
	.datac(!lpbk_lock_ack1),
	.datad(!uif_go),
	.datae(!lpbk_go),
	.dataf(!WideOr11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h002F2F2F000F0F0F;
defparam \Selector2~0 .shared_arith = "off";

dffeas \state.STATE_RMW_GO (
	.clk(mgmt_clk_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_RMW_GO~q ),
	.prn(vcc));
defparam \state.STATE_RMW_GO .is_wysiwyg = "true";
defparam \state.STATE_RMW_GO .power_up = "low";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!waitrequest_to_ctrl),
	.datab(!\state.STATE_RMW_RD~q ),
	.datac(!\state.STATE_RMW_GO~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \Selector3~0 .shared_arith = "off";

dffeas \state.STATE_RMW_RD (
	.clk(mgmt_clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_RMW_RD~q ),
	.prn(vcc));
defparam \state.STATE_RMW_RD .is_wysiwyg = "true";
defparam \state.STATE_RMW_RD .power_up = "low";

cyclonev_lcell_comb \next_state.STATE_RMW_WAIT~0 (
	.dataa(!waitrequest_to_ctrl),
	.datab(!illegal_phy_ch),
	.datac(!\state.STATE_RMW_RD~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\next_state.STATE_RMW_WAIT~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \next_state.STATE_RMW_WAIT~0 .extended_lut = "off";
defparam \next_state.STATE_RMW_WAIT~0 .lut_mask = 64'h0808080808080808;
defparam \next_state.STATE_RMW_WAIT~0 .shared_arith = "off";

dffeas \state.STATE_RMW_WAIT (
	.clk(mgmt_clk_clk),
	.d(\next_state.STATE_RMW_WAIT~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_RMW_WAIT~q ),
	.prn(vcc));
defparam \state.STATE_RMW_WAIT .is_wysiwyg = "true";
defparam \state.STATE_RMW_WAIT .power_up = "low";

dffeas \state.STATE_RMW_GO2 (
	.clk(mgmt_clk_clk),
	.d(\state.STATE_RMW_WAIT~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_RMW_GO2~q ),
	.prn(vcc));
defparam \state.STATE_RMW_GO2 .is_wysiwyg = "true";
defparam \state.STATE_RMW_GO2 .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!waitrequest_to_ctrl),
	.datab(!\state.STATE_RMW_WR~q ),
	.datac(!\state.STATE_RMW_GO2~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \Selector4~0 .shared_arith = "off";

dffeas \state.STATE_RMW_WR (
	.clk(mgmt_clk_clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_RMW_WR~q ),
	.prn(vcc));
defparam \state.STATE_RMW_WR .is_wysiwyg = "true";
defparam \state.STATE_RMW_WR .power_up = "low";

cyclonev_lcell_comb \next_state.STATE_LOCK_CHK~0 (
	.dataa(!waitrequest_to_ctrl),
	.datab(!\state.STATE_RMW_WR~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\next_state.STATE_LOCK_CHK~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \next_state.STATE_LOCK_CHK~0 .extended_lut = "off";
defparam \next_state.STATE_LOCK_CHK~0 .lut_mask = 64'h2222222222222222;
defparam \next_state.STATE_LOCK_CHK~0 .shared_arith = "off";

dffeas \state.STATE_LOCK_CHK (
	.clk(mgmt_clk_clk),
	.d(\next_state.STATE_LOCK_CHK~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_LOCK_CHK~q ),
	.prn(vcc));
defparam \state.STATE_LOCK_CHK .is_wysiwyg = "true";
defparam \state.STATE_LOCK_CHK .power_up = "low";

cyclonev_lcell_comb \next_state.STATE_GO~0 (
	.dataa(!stateSTATE_IDLE),
	.datab(!Equal6),
	.datac(!uif_go),
	.datad(!lpbk_go),
	.datae(!WideOr11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\next_state.STATE_GO~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \next_state.STATE_GO~0 .extended_lut = "off";
defparam \next_state.STATE_GO~0 .lut_mask = 64'h0888000008880000;
defparam \next_state.STATE_GO~0 .shared_arith = "off";

dffeas \state.STATE_GO (
	.clk(mgmt_clk_clk),
	.d(\next_state.STATE_GO~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_GO~q ),
	.prn(vcc));
defparam \state.STATE_GO .is_wysiwyg = "true";
defparam \state.STATE_GO .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!waitrequest_to_ctrl),
	.datab(!\state.STATE_READ~q ),
	.datac(!\state.STATE_GO~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \Selector1~0 .shared_arith = "off";

dffeas \state.STATE_READ (
	.clk(mgmt_clk_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STATE_READ~q ),
	.prn(vcc));
defparam \state.STATE_READ .is_wysiwyg = "true";
defparam \state.STATE_READ .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!lpbk_lock),
	.datab(!\state.STATE_LOCK_CHK~q ),
	.datac(!waitrequest_to_ctrl),
	.datad(!\state.STATE_READ~q ),
	.datae(!illegal_phy_ch),
	.dataf(!\state.STATE_RMW_RD~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h22F222F222F2F2F2;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~1 (
	.dataa(!stateSTATE_IDLE),
	.datab(!uif_go),
	.datac(!lpbk_go),
	.datad(!WideOr11),
	.datae(!\Selector0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~1 .extended_lut = "off";
defparam \Selector0~1 .lut_mask = 64'h7F5500007F550000;
defparam \Selector0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!lpbk_lock_ack1),
	.datab(!lpbk_lock),
	.datac(!\state.STATE_LOCK_CHK~q ),
	.datad(!uif_go),
	.datae(!lpbk_go),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h5703030357030303;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode~0 (
	.dataa(!stateSTATE_IDLE),
	.datab(!uif_go),
	.datac(!lpbk_go),
	.datad(!WideOr11),
	.datae(!\Selector5~0_combout ),
	.dataf(!\Selector0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode~0 .extended_lut = "off";
defparam \ctrl_opcode~0 .lut_mask = 64'h7F55000000000000;
defparam \ctrl_opcode~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode~1 (
	.dataa(!user_reconfig_readdata_7),
	.datab(!\next_state.STATE_GO~0_combout ),
	.datac(!\ctrl_opcode~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode~1 .extended_lut = "off";
defparam \ctrl_opcode~1 .lut_mask = 64'h0101010101010101;
defparam \ctrl_opcode~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode[0]~2 (
	.dataa(!user_reconfig_readdata_7),
	.datab(!\next_state.STATE_GO~0_combout ),
	.datac(!\ctrl_opcode~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode[0]~2 .extended_lut = "off";
defparam \ctrl_opcode[0]~2 .lut_mask = 64'h0E0E0E0E0E0E0E0E;
defparam \ctrl_opcode[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode[0]~3 (
	.dataa(!\state.STATE_RMW_WAIT~q ),
	.datab(!\ctrl_opcode[0]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode[0]~3 .extended_lut = "off";
defparam \ctrl_opcode[0]~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \ctrl_opcode[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_go~0 (
	.dataa(!\state.STATE_RMW_WAIT~q ),
	.datab(!\Selector2~0_combout ),
	.datac(!\next_state.STATE_GO~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_go~0 .extended_lut = "off";
defparam \ctrl_go~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ctrl_go~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lock~0 (
	.dataa(!\state.STATE_RMW_WAIT~q ),
	.datab(!\Selector4~0_combout ),
	.datac(!\next_state.STATE_LOCK_CHK~0_combout ),
	.datad(!\next_state.STATE_RMW_WAIT~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_lock~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lock~0 .extended_lut = "off";
defparam \ctrl_lock~0 .lut_mask = 64'h8000800080008000;
defparam \ctrl_lock~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lock~1 (
	.dataa(!lpbk_lock),
	.datab(!\Selector5~0_combout ),
	.datac(!\Selector2~0_combout ),
	.datad(!\Selector3~0_combout ),
	.datae(!\ctrl_lock~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_lock~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lock~1 .extended_lut = "off";
defparam \ctrl_lock~1 .lut_mask = 64'h5FFF1FFF5FFF1FFF;
defparam \ctrl_lock~1 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_analog_rmw_av (
	rtl,
	ifsel_notdone_resync,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_1,
	readdata_for_user_2,
	readdata_for_user_0,
	readdata_for_user_3,
	readdata_for_user_1,
	Decoder3,
	Selector2,
	analog_offset_0,
	readdata_for_user_10,
	readdata_for_user_8,
	readdata_for_user_11,
	readdata_for_user_9,
	readdata_for_user_6,
	readdata_for_user_4,
	readdata_for_user_7,
	readdata_for_user_5,
	readdata_for_user_14,
	readdata_for_user_12,
	readdata_for_user_15,
	readdata_for_user_13,
	rtl1,
	rtl2,
	readdata_for_user_16,
	WideOr4,
	WideOr41,
	analog_length,
	analog_length1,
	analog_length2,
	uif_writedata_2,
	readdata_for_user_17,
	uif_writedata_3,
	readdata_for_user_18,
	readdata_for_user_19,
	uif_writedata_5,
	readdata_for_user_20,
	uif_writedata_6,
	readdata_for_user_21,
	readdata_for_user_22,
	readdata_for_user_23,
	Equal6,
	readdata_for_user_24,
	readdata_for_user_25,
	readdata_for_user_26,
	readdata_for_user_27,
	readdata_for_user_28,
	readdata_for_user_29,
	readdata_for_user_30,
	readdata_for_user_31,
	basic_reconfig_waitrequest,
	outdata_1,
	outdata_2,
	outdata_0,
	outdata_3,
	outdata_16,
	outdata_17,
	outdata_18,
	outdata_19,
	outdata_20,
	outdata_4,
	outdata_21,
	outdata_5,
	outdata_22,
	outdata_6,
	outdata_23,
	outdata_7,
	outdata_24,
	outdata_8,
	outdata_25,
	outdata_9,
	outdata_26,
	outdata_10,
	outdata_27,
	outdata_11,
	outdata_28,
	outdata_12,
	outdata_29,
	outdata_13,
	outdata_30,
	outdata_14,
	outdata_31,
	outdata_15,
	Selector6,
	Selector61,
	result_data_0,
	rtl3,
	rtl4,
	rtl5,
	rtl6,
	rtl7,
	rtl8,
	rtl9,
	rtl10,
	rtl11,
	rtl12,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	rtl;
input 	ifsel_notdone_resync;
input 	uif_addr_offset_5;
input 	uif_addr_offset_4;
input 	uif_addr_offset_1;
input 	readdata_for_user_2;
input 	readdata_for_user_0;
input 	readdata_for_user_3;
input 	readdata_for_user_1;
input 	Decoder3;
input 	Selector2;
input 	analog_offset_0;
input 	readdata_for_user_10;
input 	readdata_for_user_8;
input 	readdata_for_user_11;
input 	readdata_for_user_9;
input 	readdata_for_user_6;
input 	readdata_for_user_4;
input 	readdata_for_user_7;
input 	readdata_for_user_5;
input 	readdata_for_user_14;
input 	readdata_for_user_12;
input 	readdata_for_user_15;
input 	readdata_for_user_13;
input 	rtl1;
input 	rtl2;
input 	readdata_for_user_16;
input 	WideOr4;
input 	WideOr41;
input 	analog_length;
input 	analog_length1;
input 	analog_length2;
input 	uif_writedata_2;
input 	readdata_for_user_17;
input 	uif_writedata_3;
input 	readdata_for_user_18;
input 	readdata_for_user_19;
input 	uif_writedata_5;
input 	readdata_for_user_20;
input 	uif_writedata_6;
input 	readdata_for_user_21;
input 	readdata_for_user_22;
input 	readdata_for_user_23;
input 	Equal6;
input 	readdata_for_user_24;
input 	readdata_for_user_25;
input 	readdata_for_user_26;
input 	readdata_for_user_27;
input 	readdata_for_user_28;
input 	readdata_for_user_29;
input 	readdata_for_user_30;
input 	readdata_for_user_31;
input 	basic_reconfig_waitrequest;
output 	outdata_1;
output 	outdata_2;
output 	outdata_0;
output 	outdata_3;
output 	outdata_16;
output 	outdata_17;
output 	outdata_18;
output 	outdata_19;
output 	outdata_20;
output 	outdata_4;
output 	outdata_21;
output 	outdata_5;
output 	outdata_22;
output 	outdata_6;
output 	outdata_23;
output 	outdata_7;
output 	outdata_24;
output 	outdata_8;
output 	outdata_25;
output 	outdata_9;
output 	outdata_26;
output 	outdata_10;
output 	outdata_27;
output 	outdata_11;
output 	outdata_28;
output 	outdata_12;
output 	outdata_29;
output 	outdata_13;
output 	outdata_30;
output 	outdata_14;
output 	outdata_31;
output 	outdata_15;
input 	Selector6;
input 	Selector61;
output 	result_data_0;
input 	rtl3;
input 	rtl4;
input 	rtl5;
input 	rtl6;
input 	rtl7;
input 	rtl8;
input 	rtl9;
input 	rtl10;
input 	rtl11;
input 	rtl12;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \result_data[1]~1_combout ;
wire \always2~0_combout ;
wire \result_data[2]~2_combout ;
wire \result_data[0]~3_combout ;
wire \result_data[0]~4_combout ;
wire \result_data[3]~5_combout ;
wire \result_data[16]~6_combout ;
wire \result_data[16]~7_combout ;
wire \result_data[18]~8_combout ;
wire \result_data[20]~9_combout ;
wire \result_data[0]~10_combout ;
wire \result_data[4]~11_combout ;
wire \result_data[4]~12_combout ;
wire \result_data[5]~13_combout ;
wire \result_data[5]~14_combout ;
wire \result_data[14]~15_combout ;
wire \wd_and_rd[6]~0_combout ;
wire \result_data[6]~16_combout ;
wire \result_data[15]~17_combout ;
wire \wd_and_rd[7]~1_combout ;
wire \result_data[7]~18_combout ;
wire \result_data[8]~19_combout ;
wire \result_data[8]~20_combout ;
wire \result_data[9]~38_combout ;
wire \result_data[10]~34_combout ;
wire \result_data[11]~21_combout ;
wire \wd_and_rd[11]~2_combout ;
wire \result_data[11]~22_combout ;
wire \result_data[12]~30_combout ;
wire \result_data[12]~26_combout ;
wire \result_data[13]~23_combout ;
wire \result_data[14]~24_combout ;
wire \result_data[15]~25_combout ;


dffeas \outdata[1] (
	.clk(mgmt_clk_clk),
	.d(\result_data[1]~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_1),
	.prn(vcc));
defparam \outdata[1] .is_wysiwyg = "true";
defparam \outdata[1] .power_up = "low";

dffeas \outdata[2] (
	.clk(mgmt_clk_clk),
	.d(\result_data[2]~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_2),
	.prn(vcc));
defparam \outdata[2] .is_wysiwyg = "true";
defparam \outdata[2] .power_up = "low";

dffeas \outdata[0] (
	.clk(mgmt_clk_clk),
	.d(\result_data[0]~4_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_0),
	.prn(vcc));
defparam \outdata[0] .is_wysiwyg = "true";
defparam \outdata[0] .power_up = "low";

dffeas \outdata[3] (
	.clk(mgmt_clk_clk),
	.d(\result_data[3]~5_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_3),
	.prn(vcc));
defparam \outdata[3] .is_wysiwyg = "true";
defparam \outdata[3] .power_up = "low";

dffeas \outdata[16] (
	.clk(mgmt_clk_clk),
	.d(\result_data[16]~7_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_16),
	.prn(vcc));
defparam \outdata[16] .is_wysiwyg = "true";
defparam \outdata[16] .power_up = "low";

dffeas \outdata[17] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_17),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_17),
	.prn(vcc));
defparam \outdata[17] .is_wysiwyg = "true";
defparam \outdata[17] .power_up = "low";

dffeas \outdata[18] (
	.clk(mgmt_clk_clk),
	.d(\result_data[18]~8_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_18),
	.prn(vcc));
defparam \outdata[18] .is_wysiwyg = "true";
defparam \outdata[18] .power_up = "low";

dffeas \outdata[19] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_19),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_19),
	.prn(vcc));
defparam \outdata[19] .is_wysiwyg = "true";
defparam \outdata[19] .power_up = "low";

dffeas \outdata[20] (
	.clk(mgmt_clk_clk),
	.d(\result_data[20]~9_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_20),
	.prn(vcc));
defparam \outdata[20] .is_wysiwyg = "true";
defparam \outdata[20] .power_up = "low";

dffeas \outdata[4] (
	.clk(mgmt_clk_clk),
	.d(\result_data[4]~12_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_4),
	.prn(vcc));
defparam \outdata[4] .is_wysiwyg = "true";
defparam \outdata[4] .power_up = "low";

dffeas \outdata[21] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_21),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_21),
	.prn(vcc));
defparam \outdata[21] .is_wysiwyg = "true";
defparam \outdata[21] .power_up = "low";

dffeas \outdata[5] (
	.clk(mgmt_clk_clk),
	.d(\result_data[5]~14_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_5),
	.prn(vcc));
defparam \outdata[5] .is_wysiwyg = "true";
defparam \outdata[5] .power_up = "low";

dffeas \outdata[22] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_22),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_22),
	.prn(vcc));
defparam \outdata[22] .is_wysiwyg = "true";
defparam \outdata[22] .power_up = "low";

dffeas \outdata[6] (
	.clk(mgmt_clk_clk),
	.d(\result_data[6]~16_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_6),
	.prn(vcc));
defparam \outdata[6] .is_wysiwyg = "true";
defparam \outdata[6] .power_up = "low";

dffeas \outdata[23] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_23),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_23),
	.prn(vcc));
defparam \outdata[23] .is_wysiwyg = "true";
defparam \outdata[23] .power_up = "low";

dffeas \outdata[7] (
	.clk(mgmt_clk_clk),
	.d(\result_data[7]~18_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_7),
	.prn(vcc));
defparam \outdata[7] .is_wysiwyg = "true";
defparam \outdata[7] .power_up = "low";

dffeas \outdata[24] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_24),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_24),
	.prn(vcc));
defparam \outdata[24] .is_wysiwyg = "true";
defparam \outdata[24] .power_up = "low";

dffeas \outdata[8] (
	.clk(mgmt_clk_clk),
	.d(\result_data[8]~20_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_8),
	.prn(vcc));
defparam \outdata[8] .is_wysiwyg = "true";
defparam \outdata[8] .power_up = "low";

dffeas \outdata[25] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_25),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_25),
	.prn(vcc));
defparam \outdata[25] .is_wysiwyg = "true";
defparam \outdata[25] .power_up = "low";

dffeas \outdata[9] (
	.clk(mgmt_clk_clk),
	.d(\result_data[9]~38_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_9),
	.prn(vcc));
defparam \outdata[9] .is_wysiwyg = "true";
defparam \outdata[9] .power_up = "low";

dffeas \outdata[26] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_26),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_26),
	.prn(vcc));
defparam \outdata[26] .is_wysiwyg = "true";
defparam \outdata[26] .power_up = "low";

dffeas \outdata[10] (
	.clk(mgmt_clk_clk),
	.d(\result_data[10]~34_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_10),
	.prn(vcc));
defparam \outdata[10] .is_wysiwyg = "true";
defparam \outdata[10] .power_up = "low";

dffeas \outdata[27] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_27),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_27),
	.prn(vcc));
defparam \outdata[27] .is_wysiwyg = "true";
defparam \outdata[27] .power_up = "low";

dffeas \outdata[11] (
	.clk(mgmt_clk_clk),
	.d(\result_data[11]~22_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_11),
	.prn(vcc));
defparam \outdata[11] .is_wysiwyg = "true";
defparam \outdata[11] .power_up = "low";

dffeas \outdata[28] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_28),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_28),
	.prn(vcc));
defparam \outdata[28] .is_wysiwyg = "true";
defparam \outdata[28] .power_up = "low";

dffeas \outdata[12] (
	.clk(mgmt_clk_clk),
	.d(\result_data[12]~26_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_12),
	.prn(vcc));
defparam \outdata[12] .is_wysiwyg = "true";
defparam \outdata[12] .power_up = "low";

dffeas \outdata[29] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_29),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_29),
	.prn(vcc));
defparam \outdata[29] .is_wysiwyg = "true";
defparam \outdata[29] .power_up = "low";

dffeas \outdata[13] (
	.clk(mgmt_clk_clk),
	.d(\result_data[13]~23_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_13),
	.prn(vcc));
defparam \outdata[13] .is_wysiwyg = "true";
defparam \outdata[13] .power_up = "low";

dffeas \outdata[30] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_30),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_30),
	.prn(vcc));
defparam \outdata[30] .is_wysiwyg = "true";
defparam \outdata[30] .power_up = "low";

dffeas \outdata[14] (
	.clk(mgmt_clk_clk),
	.d(\result_data[14]~24_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_14),
	.prn(vcc));
defparam \outdata[14] .is_wysiwyg = "true";
defparam \outdata[14] .power_up = "low";

dffeas \outdata[31] (
	.clk(mgmt_clk_clk),
	.d(readdata_for_user_31),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_31),
	.prn(vcc));
defparam \outdata[31] .is_wysiwyg = "true";
defparam \outdata[31] .power_up = "low";

dffeas \outdata[15] (
	.clk(mgmt_clk_clk),
	.d(\result_data[15]~25_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(outdata_15),
	.prn(vcc));
defparam \outdata[15] .is_wysiwyg = "true";
defparam \outdata[15] .power_up = "low";

cyclonev_lcell_comb \result_data[0]~0 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_1),
	.datad(!Decoder3),
	.datae(!Selector6),
	.dataf(!Selector61),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(result_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[0]~0 .extended_lut = "off";
defparam \result_data[0]~0 .lut_mask = 64'h0000004000AA00EA;
defparam \result_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \result_data[1]~1 (
	.dataa(!readdata_for_user_1),
	.datab(!Selector2),
	.datac(!rtl1),
	.datad(!rtl2),
	.datae(!rtl),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[1]~1 .extended_lut = "off";
defparam \result_data[1]~1 .lut_mask = 64'h1555D5555555D555;
defparam \result_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!basic_reconfig_waitrequest),
	.datab(!Equal6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h2222222222222222;
defparam \always2~0 .shared_arith = "off";

cyclonev_lcell_comb \result_data[2]~2 (
	.dataa(!readdata_for_user_2),
	.datab(!rtl1),
	.datac(!rtl2),
	.datad(!rtl4),
	.datae(!rtl5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[2]~2 .extended_lut = "off";
defparam \result_data[2]~2 .lut_mask = 64'h55D515D555D515D5;
defparam \result_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \result_data[0]~3 (
	.dataa(!analog_offset_0),
	.datab(!Selector2),
	.datac(!WideOr41),
	.datad(!analog_length),
	.datae(!analog_length2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[0]~3 .extended_lut = "off";
defparam \result_data[0]~3 .lut_mask = 64'h0888888808888888;
defparam \result_data[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \result_data[0]~4 (
	.dataa(!readdata_for_user_0),
	.datab(!rtl1),
	.datac(!rtl2),
	.datad(!\result_data[0]~3_combout ),
	.datae(!result_data_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[0]~4 .extended_lut = "off";
defparam \result_data[0]~4 .lut_mask = 64'h551555D5551555D5;
defparam \result_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \result_data[3]~5 (
	.dataa(!readdata_for_user_3),
	.datab(!rtl1),
	.datac(!rtl2),
	.datad(!rtl6),
	.datae(!rtl7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[3]~5 .extended_lut = "off";
defparam \result_data[3]~5 .lut_mask = 64'h15D555D515D555D5;
defparam \result_data[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \result_data[16]~6 (
	.dataa(!rtl2),
	.datab(!analog_length),
	.datac(!uif_writedata_2),
	.datad(!uif_writedata_6),
	.datae(!rtl8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[16]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[16]~6 .extended_lut = "off";
defparam \result_data[16]~6 .lut_mask = 64'h010101AB010101AB;
defparam \result_data[16]~6 .shared_arith = "off";

cyclonev_lcell_comb \result_data[16]~7 (
	.dataa(!rtl1),
	.datab(!rtl2),
	.datac(!readdata_for_user_16),
	.datad(!rtl8),
	.datae(!\result_data[16]~6_combout ),
	.dataf(!rtl9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[16]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[16]~7 .extended_lut = "off";
defparam \result_data[16]~7 .lut_mask = 64'h0F0B5F5F0E0A5F5F;
defparam \result_data[16]~7 .shared_arith = "off";

cyclonev_lcell_comb \result_data[18]~8 (
	.dataa(!rtl1),
	.datab(!rtl2),
	.datac(!readdata_for_user_18),
	.datad(!rtl10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[18]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[18]~8 .extended_lut = "off";
defparam \result_data[18]~8 .lut_mask = 64'h0F1F0F1F0F1F0F1F;
defparam \result_data[18]~8 .shared_arith = "off";

cyclonev_lcell_comb \result_data[20]~9 (
	.dataa(!rtl1),
	.datab(!rtl2),
	.datac(!readdata_for_user_20),
	.datad(!uif_writedata_6),
	.datae(!rtl8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[20]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[20]~9 .extended_lut = "off";
defparam \result_data[20]~9 .lut_mask = 64'h0F0F0F1F0F0F0F1F;
defparam \result_data[20]~9 .shared_arith = "off";

cyclonev_lcell_comb \result_data[0]~10 (
	.dataa(!\result_data[0]~3_combout ),
	.datab(!result_data_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[0]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[0]~10 .extended_lut = "off";
defparam \result_data[0]~10 .lut_mask = 64'h1111111111111111;
defparam \result_data[0]~10 .shared_arith = "off";

cyclonev_lcell_comb \result_data[4]~11 (
	.dataa(!rtl2),
	.datab(!analog_length),
	.datac(!uif_writedata_2),
	.datad(!\result_data[0]~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[4]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[4]~11 .extended_lut = "off";
defparam \result_data[4]~11 .lut_mask = 64'h0257025702570257;
defparam \result_data[4]~11 .shared_arith = "off";

cyclonev_lcell_comb \result_data[4]~12 (
	.dataa(!readdata_for_user_4),
	.datab(!rtl1),
	.datac(!rtl2),
	.datad(!\result_data[0]~3_combout ),
	.datae(!rtl9),
	.dataf(!\result_data[4]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[4]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[4]~12 .extended_lut = "off";
defparam \result_data[4]~12 .lut_mask = 64'h55511511DDDDDDDD;
defparam \result_data[4]~12 .shared_arith = "off";

cyclonev_lcell_comb \result_data[5]~13 (
	.dataa(!rtl2),
	.datab(!analog_length),
	.datac(!uif_writedata_3),
	.datad(!rtl11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[5]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[5]~13 .extended_lut = "off";
defparam \result_data[5]~13 .lut_mask = 64'h0257025702570257;
defparam \result_data[5]~13 .shared_arith = "off";

cyclonev_lcell_comb \result_data[5]~14 (
	.dataa(!uif_addr_offset_1),
	.datab(!readdata_for_user_5),
	.datac(!rtl1),
	.datad(!analog_length),
	.datae(!\result_data[5]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[5]~14 .extended_lut = "off";
defparam \result_data[5]~14 .lut_mask = 64'h3322F3F23322F3F2;
defparam \result_data[5]~14 .shared_arith = "off";

cyclonev_lcell_comb \result_data[14]~15 (
	.dataa(!rtl2),
	.datab(!rtl4),
	.datac(!rtl10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[14]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[14]~15 .extended_lut = "off";
defparam \result_data[14]~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \result_data[14]~15 .shared_arith = "off";

cyclonev_lcell_comb \wd_and_rd[6]~0 (
	.dataa(!rtl2),
	.datab(!rtl5),
	.datac(!rtl12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wd_and_rd[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wd_and_rd[6]~0 .extended_lut = "off";
defparam \wd_and_rd[6]~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \wd_and_rd[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \result_data[6]~16 (
	.dataa(!readdata_for_user_6),
	.datab(!rtl1),
	.datac(!\result_data[14]~15_combout ),
	.datad(!\wd_and_rd[6]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[6]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[6]~16 .extended_lut = "off";
defparam \result_data[6]~16 .lut_mask = 64'h5D1D5D1D5D1D5D1D;
defparam \result_data[6]~16 .shared_arith = "off";

cyclonev_lcell_comb \result_data[15]~17 (
	.dataa(!rtl2),
	.datab(!analog_length),
	.datac(!analog_length1),
	.datad(!uif_writedata_5),
	.datae(!rtl6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[15]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[15]~17 .extended_lut = "off";
defparam \result_data[15]~17 .lut_mask = 64'h0002555700025557;
defparam \result_data[15]~17 .shared_arith = "off";

cyclonev_lcell_comb \wd_and_rd[7]~1 (
	.dataa(!uif_addr_offset_1),
	.datab(!analog_length),
	.datac(!analog_length1),
	.datad(!rtl7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wd_and_rd[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wd_and_rd[7]~1 .extended_lut = "off";
defparam \wd_and_rd[7]~1 .lut_mask = 64'h2301230123012301;
defparam \wd_and_rd[7]~1 .shared_arith = "off";

cyclonev_lcell_comb \result_data[7]~18 (
	.dataa(!readdata_for_user_7),
	.datab(!rtl1),
	.datac(!\result_data[15]~17_combout ),
	.datad(!\wd_and_rd[7]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[7]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[7]~18 .extended_lut = "off";
defparam \result_data[7]~18 .lut_mask = 64'h5D0C5D0C5D0C5D0C;
defparam \result_data[7]~18 .shared_arith = "off";

cyclonev_lcell_comb \result_data[8]~19 (
	.dataa(!uif_addr_offset_1),
	.datab(!readdata_for_user_8),
	.datac(!WideOr4),
	.datad(!analog_length),
	.datae(!analog_length1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[8]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[8]~19 .extended_lut = "off";
defparam \result_data[8]~19 .lut_mask = 64'h3311331033113310;
defparam \result_data[8]~19 .shared_arith = "off";

cyclonev_lcell_comb \result_data[8]~20 (
	.dataa(!rtl1),
	.datab(!rtl2),
	.datac(!\result_data[0]~10_combout ),
	.datad(!\result_data[16]~6_combout ),
	.datae(!\result_data[8]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[8]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[8]~20 .extended_lut = "off";
defparam \result_data[8]~20 .lut_mask = 64'h04AEFFFF04AEFFFF;
defparam \result_data[8]~20 .shared_arith = "off";

cyclonev_lcell_comb \result_data[9]~38 (
	.dataa(!readdata_for_user_9),
	.datab(!uif_addr_offset_1),
	.datac(!uif_writedata_3),
	.datad(!analog_length),
	.datae(!rtl2),
	.dataf(!rtl1),
	.datag(!rtl11),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[9]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[9]~38 .extended_lut = "on";
defparam \result_data[9]~38 .lut_mask = 64'h5511551F5F1F5511;
defparam \result_data[9]~38 .shared_arith = "off";

cyclonev_lcell_comb \result_data[10]~34 (
	.dataa(!rtl12),
	.datab(!rtl5),
	.datac(!rtl10),
	.datad(!readdata_for_user_10),
	.datae(!rtl2),
	.dataf(!rtl1),
	.datag(!rtl4),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[10]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[10]~34 .extended_lut = "on";
defparam \result_data[10]~34 .lut_mask = 64'h00FF0FAF0FCF00FF;
defparam \result_data[10]~34 .shared_arith = "off";

cyclonev_lcell_comb \result_data[11]~21 (
	.dataa(!rtl1),
	.datab(!analog_length),
	.datac(!analog_length1),
	.datad(!uif_writedata_5),
	.datae(!rtl6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[11]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[11]~21 .extended_lut = "off";
defparam \result_data[11]~21 .lut_mask = 64'h0002555700025557;
defparam \result_data[11]~21 .shared_arith = "off";

cyclonev_lcell_comb \wd_and_rd[11]~2 (
	.dataa(!analog_offset_0),
	.datab(!Selector2),
	.datac(!analog_length),
	.datad(!analog_length2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wd_and_rd[11]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wd_and_rd[11]~2 .extended_lut = "off";
defparam \wd_and_rd[11]~2 .lut_mask = 64'h0002000200020002;
defparam \wd_and_rd[11]~2 .shared_arith = "off";

cyclonev_lcell_comb \result_data[11]~22 (
	.dataa(!readdata_for_user_11),
	.datab(!rtl1),
	.datac(!rtl2),
	.datad(!rtl7),
	.datae(!\result_data[11]~21_combout ),
	.dataf(!\wd_and_rd[11]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[11]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[11]~22 .extended_lut = "off";
defparam \result_data[11]~22 .lut_mask = 64'h45557D7D41517D7D;
defparam \result_data[11]~22 .shared_arith = "off";

cyclonev_lcell_comb \result_data[12]~30 (
	.dataa(!uif_writedata_2),
	.datab(!analog_length),
	.datac(!result_data_0),
	.datad(!rtl2),
	.datae(!\result_data[0]~3_combout ),
	.dataf(!rtl1),
	.datag(!readdata_for_user_12),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[12]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[12]~30 .extended_lut = "on";
defparam \result_data[12]~30 .lut_mask = 64'h00000000110F110F;
defparam \result_data[12]~30 .shared_arith = "off";

cyclonev_lcell_comb \result_data[12]~26 (
	.dataa(!rtl8),
	.datab(!\result_data[12]~30_combout ),
	.datac(!rtl9),
	.datad(!rtl2),
	.datae(!rtl1),
	.dataf(!readdata_for_user_12),
	.datag(!uif_writedata_6),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[12]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[12]~26 .extended_lut = "on";
defparam \result_data[12]~26 .lut_mask = 64'h33373333FFBFF333;
defparam \result_data[12]~26 .shared_arith = "off";

cyclonev_lcell_comb \result_data[13]~23 (
	.dataa(!readdata_for_user_13),
	.datab(!rtl1),
	.datac(!\result_data[5]~13_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[13]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[13]~23 .extended_lut = "off";
defparam \result_data[13]~23 .lut_mask = 64'h5757575757575757;
defparam \result_data[13]~23 .shared_arith = "off";

cyclonev_lcell_comb \result_data[14]~24 (
	.dataa(!readdata_for_user_14),
	.datab(!rtl1),
	.datac(!\result_data[14]~15_combout ),
	.datad(!\wd_and_rd[6]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[14]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[14]~24 .extended_lut = "off";
defparam \result_data[14]~24 .lut_mask = 64'h5747574757475747;
defparam \result_data[14]~24 .shared_arith = "off";

cyclonev_lcell_comb \result_data[15]~25 (
	.dataa(!readdata_for_user_15),
	.datab(!rtl1),
	.datac(!rtl2),
	.datad(!rtl7),
	.datae(!\result_data[15]~17_combout ),
	.dataf(!\wd_and_rd[11]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\result_data[15]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_data[15]~25 .extended_lut = "off";
defparam \result_data[15]~25 .lut_mask = 64'h5455777744457777;
defparam \result_data[15]~25 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_cif (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_11,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write,
	grant_1,
	mutex_req,
	master_address_2,
	mutex_grant,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	ifsel_notdone_resync,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_0,
	uif_addr_offset_1,
	uif_addr_offset_3,
	readdata_for_user_2,
	readdata_for_user_0,
	readdata_for_user_3,
	readdata_for_user_1,
	Decoder3,
	lpbk_lock,
	readdata_for_user_10,
	readdata_for_user_8,
	readdata_for_user_11,
	readdata_for_user_9,
	readdata_for_user_6,
	readdata_for_user_4,
	readdata_for_user_7,
	readdata_for_user_5,
	readdata_for_user_14,
	readdata_for_user_12,
	readdata_for_user_15,
	readdata_for_user_13,
	readdata_for_user_16,
	analog_length,
	uif_logical_ch_addr_0,
	ph_readdata_0,
	uif_logical_ch_addr_1,
	ph_readdata_1,
	readdata_for_user_17,
	uif_logical_ch_addr_2,
	ph_readdata_2,
	readdata_for_user_18,
	uif_logical_ch_addr_3,
	ph_readdata_3,
	readdata_for_user_19,
	uif_logical_ch_addr_4,
	ph_readdata_4,
	readdata_for_user_20,
	uif_logical_ch_addr_5,
	ph_readdata_5,
	readdata_for_user_21,
	ph_readdata_6,
	uif_logical_ch_addr_6,
	readdata_for_user_22,
	ph_readdata_7,
	uif_logical_ch_addr_7,
	readdata_for_user_23,
	uif_logical_ch_addr_8,
	ph_readdata_8,
	readdata_for_user_24,
	ph_readdata_9,
	uif_logical_ch_addr_9,
	ph_readdata_10,
	readdata_for_user_25,
	ph_readdata_11,
	readdata_for_user_26,
	ph_readdata_12,
	readdata_for_user_27,
	ph_readdata_13,
	readdata_for_user_28,
	ph_readdata_14,
	readdata_for_user_29,
	ph_readdata_15,
	readdata_for_user_30,
	ph_readdata_16,
	readdata_for_user_31,
	ph_readdata_17,
	ph_readdata_18,
	ph_readdata_19,
	ph_readdata_20,
	ph_readdata_21,
	ph_readdata_22,
	ph_readdata_23,
	ph_readdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	ctrl_opcode_1,
	ctrl_opcode_0,
	ctrl_go,
	ctrl_lock,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	waitrequest_to_ctrl,
	illegal_phy_ch,
	outdata_1,
	outdata_2,
	outdata_0,
	outdata_3,
	outdata_16,
	outdata_17,
	outdata_18,
	outdata_19,
	outdata_20,
	WideOr5,
	outdata_4,
	outdata_21,
	outdata_5,
	outdata_22,
	outdata_6,
	outdata_23,
	outdata_7,
	outdata_24,
	outdata_8,
	outdata_25,
	outdata_9,
	outdata_26,
	outdata_10,
	outdata_27,
	outdata_11,
	outdata_28,
	outdata_12,
	outdata_29,
	outdata_13,
	outdata_30,
	outdata_14,
	outdata_31,
	outdata_15,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_16;
input 	basic_reconfig_readdata_17;
input 	basic_reconfig_readdata_18;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	master_writedata_16;
output 	master_writedata_17;
output 	master_writedata_18;
output 	master_writedata_19;
output 	master_writedata_20;
output 	master_writedata_21;
output 	master_writedata_22;
output 	master_writedata_23;
output 	master_writedata_24;
output 	master_writedata_25;
output 	master_writedata_26;
output 	master_writedata_27;
output 	master_writedata_11;
output 	master_writedata_28;
output 	master_writedata_12;
output 	master_writedata_29;
output 	master_writedata_13;
output 	master_writedata_30;
output 	master_writedata_14;
output 	master_writedata_31;
output 	master_writedata_15;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write;
input 	grant_1;
output 	mutex_req;
output 	master_address_2;
output 	mutex_grant;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	ifsel_notdone_resync;
input 	uif_addr_offset_5;
input 	uif_addr_offset_4;
input 	uif_addr_offset_0;
input 	uif_addr_offset_1;
input 	uif_addr_offset_3;
output 	readdata_for_user_2;
output 	readdata_for_user_0;
output 	readdata_for_user_3;
output 	readdata_for_user_1;
input 	Decoder3;
input 	lpbk_lock;
output 	readdata_for_user_10;
output 	readdata_for_user_8;
output 	readdata_for_user_11;
output 	readdata_for_user_9;
output 	readdata_for_user_6;
output 	readdata_for_user_4;
output 	readdata_for_user_7;
output 	readdata_for_user_5;
output 	readdata_for_user_14;
output 	readdata_for_user_12;
output 	readdata_for_user_15;
output 	readdata_for_user_13;
output 	readdata_for_user_16;
input 	analog_length;
input 	uif_logical_ch_addr_0;
output 	ph_readdata_0;
input 	uif_logical_ch_addr_1;
output 	ph_readdata_1;
output 	readdata_for_user_17;
input 	uif_logical_ch_addr_2;
output 	ph_readdata_2;
output 	readdata_for_user_18;
input 	uif_logical_ch_addr_3;
output 	ph_readdata_3;
output 	readdata_for_user_19;
input 	uif_logical_ch_addr_4;
output 	ph_readdata_4;
output 	readdata_for_user_20;
input 	uif_logical_ch_addr_5;
output 	ph_readdata_5;
output 	readdata_for_user_21;
output 	ph_readdata_6;
input 	uif_logical_ch_addr_6;
output 	readdata_for_user_22;
output 	ph_readdata_7;
input 	uif_logical_ch_addr_7;
output 	readdata_for_user_23;
input 	uif_logical_ch_addr_8;
output 	ph_readdata_8;
output 	readdata_for_user_24;
output 	ph_readdata_9;
input 	uif_logical_ch_addr_9;
output 	ph_readdata_10;
output 	readdata_for_user_25;
output 	ph_readdata_11;
output 	readdata_for_user_26;
output 	ph_readdata_12;
output 	readdata_for_user_27;
output 	ph_readdata_13;
output 	readdata_for_user_28;
output 	ph_readdata_14;
output 	readdata_for_user_29;
output 	ph_readdata_15;
output 	readdata_for_user_30;
output 	ph_readdata_16;
output 	readdata_for_user_31;
output 	ph_readdata_17;
output 	ph_readdata_18;
output 	ph_readdata_19;
output 	ph_readdata_20;
output 	ph_readdata_21;
output 	ph_readdata_22;
output 	ph_readdata_23;
output 	ph_readdata_24;
output 	ph_readdata_25;
output 	ph_readdata_26;
output 	ph_readdata_27;
output 	ph_readdata_28;
output 	ph_readdata_29;
output 	ph_readdata_30;
output 	ph_readdata_31;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	ctrl_opcode_1;
input 	ctrl_opcode_0;
input 	ctrl_go;
input 	ctrl_lock;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	waitrequest_to_ctrl;
output 	illegal_phy_ch;
input 	outdata_1;
input 	outdata_2;
input 	outdata_0;
input 	outdata_3;
input 	outdata_16;
input 	outdata_17;
input 	outdata_18;
input 	outdata_19;
input 	outdata_20;
input 	WideOr5;
input 	outdata_4;
input 	outdata_21;
input 	outdata_5;
input 	outdata_22;
input 	outdata_6;
input 	outdata_23;
input 	outdata_7;
input 	outdata_24;
input 	outdata_8;
input 	outdata_25;
input 	outdata_9;
input 	outdata_26;
input 	outdata_10;
input 	outdata_27;
input 	outdata_11;
input 	outdata_28;
input 	outdata_12;
input 	outdata_29;
input 	outdata_13;
input 	outdata_30;
input 	outdata_14;
input 	outdata_31;
input 	outdata_15;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



RECONFIGURE_IP_alt_arbiter_acq mutex_inst(
	.grant_1(grant_1),
	.mutex_req(mutex_req),
	.mutex_grant1(mutex_grant));

RECONFIGURE_IP_alt_xreconf_basic_acq inst_basic_acq(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.master_writedata_16(master_writedata_16),
	.master_writedata_17(master_writedata_17),
	.master_writedata_18(master_writedata_18),
	.master_writedata_19(master_writedata_19),
	.master_writedata_20(master_writedata_20),
	.master_writedata_21(master_writedata_21),
	.master_writedata_22(master_writedata_22),
	.master_writedata_23(master_writedata_23),
	.master_writedata_24(master_writedata_24),
	.master_writedata_25(master_writedata_25),
	.master_writedata_26(master_writedata_26),
	.master_writedata_27(master_writedata_27),
	.master_writedata_11(master_writedata_11),
	.master_writedata_28(master_writedata_28),
	.master_writedata_12(master_writedata_12),
	.master_writedata_29(master_writedata_29),
	.master_writedata_13(master_writedata_13),
	.master_writedata_30(master_writedata_30),
	.master_writedata_14(master_writedata_14),
	.master_writedata_31(master_writedata_31),
	.master_writedata_15(master_writedata_15),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.master_write1(master_write),
	.mutex_req1(mutex_req),
	.master_address_2(master_address_2),
	.mutex_grant(mutex_grant),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read1(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.reset(ifsel_notdone_resync),
	.uif_addr_offset_5(uif_addr_offset_5),
	.uif_addr_offset_4(uif_addr_offset_4),
	.uif_addr_offset_0(uif_addr_offset_0),
	.uif_addr_offset_1(uif_addr_offset_1),
	.uif_addr_offset_3(uif_addr_offset_3),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_1(readdata_for_user_1),
	.Decoder3(Decoder3),
	.lpbk_lock(lpbk_lock),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_9(readdata_for_user_9),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_13(readdata_for_user_13),
	.readdata_for_user_16(readdata_for_user_16),
	.analog_length(analog_length),
	.logical_ch_addr({uif_logical_ch_addr_9,uif_logical_ch_addr_8,uif_logical_ch_addr_7,uif_logical_ch_addr_6,uif_logical_ch_addr_5,uif_logical_ch_addr_4,uif_logical_ch_addr_3,uif_logical_ch_addr_2,uif_logical_ch_addr_1,uif_logical_ch_addr_0}),
	.ph_readdata_0(ph_readdata_0),
	.ph_readdata_1(ph_readdata_1),
	.readdata_for_user_17(readdata_for_user_17),
	.ph_readdata_2(ph_readdata_2),
	.readdata_for_user_18(readdata_for_user_18),
	.ph_readdata_3(ph_readdata_3),
	.readdata_for_user_19(readdata_for_user_19),
	.ph_readdata_4(ph_readdata_4),
	.readdata_for_user_20(readdata_for_user_20),
	.ph_readdata_5(ph_readdata_5),
	.readdata_for_user_21(readdata_for_user_21),
	.ph_readdata_6(ph_readdata_6),
	.readdata_for_user_22(readdata_for_user_22),
	.ph_readdata_7(ph_readdata_7),
	.readdata_for_user_23(readdata_for_user_23),
	.ph_readdata_8(ph_readdata_8),
	.readdata_for_user_24(readdata_for_user_24),
	.ph_readdata_9(ph_readdata_9),
	.ph_readdata_10(ph_readdata_10),
	.readdata_for_user_25(readdata_for_user_25),
	.ph_readdata_11(ph_readdata_11),
	.readdata_for_user_26(readdata_for_user_26),
	.ph_readdata_12(ph_readdata_12),
	.readdata_for_user_27(readdata_for_user_27),
	.ph_readdata_13(ph_readdata_13),
	.readdata_for_user_28(readdata_for_user_28),
	.ph_readdata_14(ph_readdata_14),
	.readdata_for_user_29(readdata_for_user_29),
	.ph_readdata_15(ph_readdata_15),
	.readdata_for_user_30(readdata_for_user_30),
	.ph_readdata_16(ph_readdata_16),
	.readdata_for_user_31(readdata_for_user_31),
	.ph_readdata_17(ph_readdata_17),
	.ph_readdata_18(ph_readdata_18),
	.ph_readdata_19(ph_readdata_19),
	.ph_readdata_20(ph_readdata_20),
	.ph_readdata_21(ph_readdata_21),
	.ph_readdata_22(ph_readdata_22),
	.ph_readdata_23(ph_readdata_23),
	.ph_readdata_24(ph_readdata_24),
	.ph_readdata_25(ph_readdata_25),
	.ph_readdata_26(ph_readdata_26),
	.ph_readdata_27(ph_readdata_27),
	.ph_readdata_28(ph_readdata_28),
	.ph_readdata_29(ph_readdata_29),
	.ph_readdata_30(ph_readdata_30),
	.ph_readdata_31(ph_readdata_31),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.ctrl_opcode_1(ctrl_opcode_1),
	.ctrl_opcode_0(ctrl_opcode_0),
	.ctrl_go(ctrl_go),
	.ctrl_lock(ctrl_lock),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.waitrequest_to_ctrl1(waitrequest_to_ctrl),
	.illegal_phy_ch1(illegal_phy_ch),
	.outdata_1(outdata_1),
	.outdata_2(outdata_2),
	.outdata_0(outdata_0),
	.outdata_3(outdata_3),
	.outdata_16(outdata_16),
	.outdata_17(outdata_17),
	.outdata_18(outdata_18),
	.outdata_19(outdata_19),
	.outdata_20(outdata_20),
	.WideOr5(WideOr5),
	.outdata_4(outdata_4),
	.outdata_21(outdata_21),
	.outdata_5(outdata_5),
	.outdata_22(outdata_22),
	.outdata_6(outdata_6),
	.outdata_23(outdata_23),
	.outdata_7(outdata_7),
	.outdata_24(outdata_24),
	.outdata_8(outdata_8),
	.outdata_25(outdata_25),
	.outdata_9(outdata_9),
	.outdata_26(outdata_26),
	.outdata_10(outdata_10),
	.outdata_27(outdata_27),
	.outdata_11(outdata_11),
	.outdata_28(outdata_28),
	.outdata_12(outdata_12),
	.outdata_29(outdata_29),
	.outdata_13(outdata_13),
	.outdata_30(outdata_30),
	.outdata_14(outdata_14),
	.outdata_31(outdata_31),
	.outdata_15(outdata_15),
	.clk(mgmt_clk_clk));

endmodule

module RECONFIGURE_IP_alt_arbiter_acq (
	grant_1,
	mutex_req,
	mutex_grant1)/* synthesis synthesis_greybox=0 */;
input 	grant_1;
input 	mutex_req;
output 	mutex_grant1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb mutex_grant(
	.dataa(!grant_1),
	.datab(!mutex_req),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mutex_grant1),
	.sumout(),
	.cout(),
	.shareout());
defparam mutex_grant.extended_lut = "off";
defparam mutex_grant.lut_mask = 64'h1111111111111111;
defparam mutex_grant.shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_basic_acq (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_11,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write1,
	mutex_req1,
	master_address_2,
	mutex_grant,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read1,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	reset,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_0,
	uif_addr_offset_1,
	uif_addr_offset_3,
	readdata_for_user_2,
	readdata_for_user_0,
	readdata_for_user_3,
	readdata_for_user_1,
	Decoder3,
	lpbk_lock,
	readdata_for_user_10,
	readdata_for_user_8,
	readdata_for_user_11,
	readdata_for_user_9,
	readdata_for_user_6,
	readdata_for_user_4,
	readdata_for_user_7,
	readdata_for_user_5,
	readdata_for_user_14,
	readdata_for_user_12,
	readdata_for_user_15,
	readdata_for_user_13,
	readdata_for_user_16,
	analog_length,
	logical_ch_addr,
	ph_readdata_0,
	ph_readdata_1,
	readdata_for_user_17,
	ph_readdata_2,
	readdata_for_user_18,
	ph_readdata_3,
	readdata_for_user_19,
	ph_readdata_4,
	readdata_for_user_20,
	ph_readdata_5,
	readdata_for_user_21,
	ph_readdata_6,
	readdata_for_user_22,
	ph_readdata_7,
	readdata_for_user_23,
	ph_readdata_8,
	readdata_for_user_24,
	ph_readdata_9,
	ph_readdata_10,
	readdata_for_user_25,
	ph_readdata_11,
	readdata_for_user_26,
	ph_readdata_12,
	readdata_for_user_27,
	ph_readdata_13,
	readdata_for_user_28,
	ph_readdata_14,
	readdata_for_user_29,
	ph_readdata_15,
	readdata_for_user_30,
	ph_readdata_16,
	readdata_for_user_31,
	ph_readdata_17,
	ph_readdata_18,
	ph_readdata_19,
	ph_readdata_20,
	ph_readdata_21,
	ph_readdata_22,
	ph_readdata_23,
	ph_readdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	ctrl_opcode_1,
	ctrl_opcode_0,
	ctrl_go,
	ctrl_lock,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	waitrequest_to_ctrl1,
	illegal_phy_ch1,
	outdata_1,
	outdata_2,
	outdata_0,
	outdata_3,
	outdata_16,
	outdata_17,
	outdata_18,
	outdata_19,
	outdata_20,
	WideOr5,
	outdata_4,
	outdata_21,
	outdata_5,
	outdata_22,
	outdata_6,
	outdata_23,
	outdata_7,
	outdata_24,
	outdata_8,
	outdata_25,
	outdata_9,
	outdata_26,
	outdata_10,
	outdata_27,
	outdata_11,
	outdata_28,
	outdata_12,
	outdata_29,
	outdata_13,
	outdata_30,
	outdata_14,
	outdata_31,
	outdata_15,
	clk)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_16;
input 	basic_reconfig_readdata_17;
input 	basic_reconfig_readdata_18;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	master_writedata_16;
output 	master_writedata_17;
output 	master_writedata_18;
output 	master_writedata_19;
output 	master_writedata_20;
output 	master_writedata_21;
output 	master_writedata_22;
output 	master_writedata_23;
output 	master_writedata_24;
output 	master_writedata_25;
output 	master_writedata_26;
output 	master_writedata_27;
output 	master_writedata_11;
output 	master_writedata_28;
output 	master_writedata_12;
output 	master_writedata_29;
output 	master_writedata_13;
output 	master_writedata_30;
output 	master_writedata_14;
output 	master_writedata_31;
output 	master_writedata_15;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write1;
output 	mutex_req1;
output 	master_address_2;
input 	mutex_grant;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read1;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	reset;
input 	uif_addr_offset_5;
input 	uif_addr_offset_4;
input 	uif_addr_offset_0;
input 	uif_addr_offset_1;
input 	uif_addr_offset_3;
output 	readdata_for_user_2;
output 	readdata_for_user_0;
output 	readdata_for_user_3;
output 	readdata_for_user_1;
input 	Decoder3;
input 	lpbk_lock;
output 	readdata_for_user_10;
output 	readdata_for_user_8;
output 	readdata_for_user_11;
output 	readdata_for_user_9;
output 	readdata_for_user_6;
output 	readdata_for_user_4;
output 	readdata_for_user_7;
output 	readdata_for_user_5;
output 	readdata_for_user_14;
output 	readdata_for_user_12;
output 	readdata_for_user_15;
output 	readdata_for_user_13;
output 	readdata_for_user_16;
input 	analog_length;
input 	[9:0] logical_ch_addr;
output 	ph_readdata_0;
output 	ph_readdata_1;
output 	readdata_for_user_17;
output 	ph_readdata_2;
output 	readdata_for_user_18;
output 	ph_readdata_3;
output 	readdata_for_user_19;
output 	ph_readdata_4;
output 	readdata_for_user_20;
output 	ph_readdata_5;
output 	readdata_for_user_21;
output 	ph_readdata_6;
output 	readdata_for_user_22;
output 	ph_readdata_7;
output 	readdata_for_user_23;
output 	ph_readdata_8;
output 	readdata_for_user_24;
output 	ph_readdata_9;
output 	ph_readdata_10;
output 	readdata_for_user_25;
output 	ph_readdata_11;
output 	readdata_for_user_26;
output 	ph_readdata_12;
output 	readdata_for_user_27;
output 	ph_readdata_13;
output 	readdata_for_user_28;
output 	ph_readdata_14;
output 	readdata_for_user_29;
output 	ph_readdata_15;
output 	readdata_for_user_30;
output 	ph_readdata_16;
output 	readdata_for_user_31;
output 	ph_readdata_17;
output 	ph_readdata_18;
output 	ph_readdata_19;
output 	ph_readdata_20;
output 	ph_readdata_21;
output 	ph_readdata_22;
output 	ph_readdata_23;
output 	ph_readdata_24;
output 	ph_readdata_25;
output 	ph_readdata_26;
output 	ph_readdata_27;
output 	ph_readdata_28;
output 	ph_readdata_29;
output 	ph_readdata_30;
output 	ph_readdata_31;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	ctrl_opcode_1;
input 	ctrl_opcode_0;
input 	ctrl_go;
input 	ctrl_lock;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	waitrequest_to_ctrl1;
output 	illegal_phy_ch1;
input 	outdata_1;
input 	outdata_2;
input 	outdata_0;
input 	outdata_3;
input 	outdata_16;
input 	outdata_17;
input 	outdata_18;
input 	outdata_19;
input 	outdata_20;
input 	WideOr5;
input 	outdata_4;
input 	outdata_21;
input 	outdata_5;
input 	outdata_22;
input 	outdata_6;
input 	outdata_23;
input 	outdata_7;
input 	outdata_24;
input 	outdata_8;
input 	outdata_25;
input 	outdata_9;
input 	outdata_26;
input 	outdata_10;
input 	outdata_27;
input 	outdata_11;
input 	outdata_28;
input 	outdata_12;
input 	outdata_29;
input 	outdata_13;
input 	outdata_30;
input 	outdata_14;
input 	outdata_31;
input 	outdata_15;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lch_dly[7]~q ;
wire \lch_dly[5]~q ;
wire \lch_dly[6]~q ;
wire \lch_legal~0_combout ;
wire \lch_dly[8]~q ;
wire \lch_dly[9]~q ;
wire \lch_legal~1_combout ;
wire \lch_dly[4]~q ;
wire \Selector5~2_combout ;
wire \lch_dly[0]~q ;
wire \lch_dly[1]~q ;
wire \lch_legal~2_combout ;
wire \lch_dly[2]~q ;
wire \lch_dly[3]~q ;
wire \lch_legal~3_combout ;
wire \lch_legal~4_combout ;
wire \lch_legal~5_combout ;
wire \lch_legal~6_combout ;
wire \lch_legal~q ;
wire \state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ;
wire \Selector9~0_combout ;
wire \state.ST_SET_RECONFIG_BASIC_WRITE~q ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ;
wire \Selector13~0_combout ;
wire \state.ST_START_AGAIN~q ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ;
wire \Selector5~4_combout ;
wire \Selector5~5_combout ;
wire \Selector5~6_combout ;
wire \Selector5~7_combout ;
wire \Selector10~0_combout ;
wire \state.ST_SET_RECONFIG_BASIC_READ~q ;
wire \Selector11~0_combout ;
wire \state.ST_READ_RECONFIG_BASIC_DATA~q ;
wire \Selector12~0_combout ;
wire \Selector12~1_combout ;
wire \state.ST_CHECK_CTRLLOCK~q ;
wire \Selector14~0_combout ;
wire \state.ST_RELEASE_REQ~q ;
wire \Selector0~0_combout ;
wire \state.0000~q ;
wire \Selector1~0_combout ;
wire \state.ST_REQ_MUTEX~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \state.ST_WRITE_RECONFIG_BASIC_LCH~q ;
wire \Selector3~0_combout ;
wire \state.ST_READ_PHY_ADDRESS~q ;
wire \Selector4~0_combout ;
wire \state.ST_CHECK_PHY_ADD_LEGAL~q ;
wire \Selector5~3_combout ;
wire \Selector8~0_combout ;
wire \WideOr7~0_combout ;
wire \WideOr8~combout ;
wire \WideOr5~0_combout ;
wire \WideOr17~0_combout ;
wire \Selector28~0_combout ;
wire \WideOr7~combout ;
wire \WideOr6~combout ;
wire \WideOr9~combout ;
wire \Selector12~2_combout ;
wire \readdata_for_user[0]~0_combout ;
wire \Selector16~0_combout ;
wire \ph_readdata[6]~0_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \Selector25~0_combout ;
wire \Selector25~1_combout ;
wire \Selector27~0_combout ;
wire \Selector27~1_combout ;
wire \Selector27~2_combout ;
wire \Selector24~0_combout ;
wire \Selector24~1_combout ;
wire \Selector23~0_combout ;
wire \Selector23~1_combout ;
wire \Selector22~0_combout ;
wire \Selector21~0_combout ;
wire \Selector20~0_combout ;
wire \Selector19~0_combout ;
wire \Selector18~0_combout ;
wire \Selector17~0_combout ;
wire \Selector16~1_combout ;


dffeas \master_writedata[16] (
	.clk(clk),
	.d(outdata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_16),
	.prn(vcc));
defparam \master_writedata[16] .is_wysiwyg = "true";
defparam \master_writedata[16] .power_up = "low";

dffeas \master_writedata[17] (
	.clk(clk),
	.d(outdata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_17),
	.prn(vcc));
defparam \master_writedata[17] .is_wysiwyg = "true";
defparam \master_writedata[17] .power_up = "low";

dffeas \master_writedata[18] (
	.clk(clk),
	.d(outdata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_18),
	.prn(vcc));
defparam \master_writedata[18] .is_wysiwyg = "true";
defparam \master_writedata[18] .power_up = "low";

dffeas \master_writedata[19] (
	.clk(clk),
	.d(outdata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_19),
	.prn(vcc));
defparam \master_writedata[19] .is_wysiwyg = "true";
defparam \master_writedata[19] .power_up = "low";

dffeas \master_writedata[20] (
	.clk(clk),
	.d(outdata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_20),
	.prn(vcc));
defparam \master_writedata[20] .is_wysiwyg = "true";
defparam \master_writedata[20] .power_up = "low";

dffeas \master_writedata[21] (
	.clk(clk),
	.d(outdata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_21),
	.prn(vcc));
defparam \master_writedata[21] .is_wysiwyg = "true";
defparam \master_writedata[21] .power_up = "low";

dffeas \master_writedata[22] (
	.clk(clk),
	.d(outdata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_22),
	.prn(vcc));
defparam \master_writedata[22] .is_wysiwyg = "true";
defparam \master_writedata[22] .power_up = "low";

dffeas \master_writedata[23] (
	.clk(clk),
	.d(outdata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_23),
	.prn(vcc));
defparam \master_writedata[23] .is_wysiwyg = "true";
defparam \master_writedata[23] .power_up = "low";

dffeas \master_writedata[24] (
	.clk(clk),
	.d(outdata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_24),
	.prn(vcc));
defparam \master_writedata[24] .is_wysiwyg = "true";
defparam \master_writedata[24] .power_up = "low";

dffeas \master_writedata[25] (
	.clk(clk),
	.d(outdata_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_25),
	.prn(vcc));
defparam \master_writedata[25] .is_wysiwyg = "true";
defparam \master_writedata[25] .power_up = "low";

dffeas \master_writedata[26] (
	.clk(clk),
	.d(outdata_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_26),
	.prn(vcc));
defparam \master_writedata[26] .is_wysiwyg = "true";
defparam \master_writedata[26] .power_up = "low";

dffeas \master_writedata[27] (
	.clk(clk),
	.d(outdata_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_27),
	.prn(vcc));
defparam \master_writedata[27] .is_wysiwyg = "true";
defparam \master_writedata[27] .power_up = "low";

dffeas \master_writedata[11] (
	.clk(clk),
	.d(outdata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_11),
	.prn(vcc));
defparam \master_writedata[11] .is_wysiwyg = "true";
defparam \master_writedata[11] .power_up = "low";

dffeas \master_writedata[28] (
	.clk(clk),
	.d(outdata_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_28),
	.prn(vcc));
defparam \master_writedata[28] .is_wysiwyg = "true";
defparam \master_writedata[28] .power_up = "low";

dffeas \master_writedata[12] (
	.clk(clk),
	.d(outdata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_12),
	.prn(vcc));
defparam \master_writedata[12] .is_wysiwyg = "true";
defparam \master_writedata[12] .power_up = "low";

dffeas \master_writedata[29] (
	.clk(clk),
	.d(outdata_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_29),
	.prn(vcc));
defparam \master_writedata[29] .is_wysiwyg = "true";
defparam \master_writedata[29] .power_up = "low";

dffeas \master_writedata[13] (
	.clk(clk),
	.d(outdata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_13),
	.prn(vcc));
defparam \master_writedata[13] .is_wysiwyg = "true";
defparam \master_writedata[13] .power_up = "low";

dffeas \master_writedata[30] (
	.clk(clk),
	.d(outdata_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_30),
	.prn(vcc));
defparam \master_writedata[30] .is_wysiwyg = "true";
defparam \master_writedata[30] .power_up = "low";

dffeas \master_writedata[14] (
	.clk(clk),
	.d(outdata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_14),
	.prn(vcc));
defparam \master_writedata[14] .is_wysiwyg = "true";
defparam \master_writedata[14] .power_up = "low";

dffeas \master_writedata[31] (
	.clk(clk),
	.d(outdata_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_31),
	.prn(vcc));
defparam \master_writedata[31] .is_wysiwyg = "true";
defparam \master_writedata[31] .power_up = "low";

dffeas \master_writedata[15] (
	.clk(clk),
	.d(outdata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!\Selector8~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_15),
	.prn(vcc));
defparam \master_writedata[15] .is_wysiwyg = "true";
defparam \master_writedata[15] .power_up = "low";

dffeas master_write(
	.clk(clk),
	.d(\WideOr8~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write1),
	.prn(vcc));
defparam master_write.is_wysiwyg = "true";
defparam master_write.power_up = "low";

dffeas mutex_req(
	.clk(clk),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mutex_req1),
	.prn(vcc));
defparam mutex_req.is_wysiwyg = "true";
defparam mutex_req.power_up = "low";

dffeas \master_address[2] (
	.clk(clk),
	.d(\WideOr5~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_2),
	.prn(vcc));
defparam \master_address[2] .is_wysiwyg = "true";
defparam \master_address[2] .power_up = "low";

dffeas \master_address[0] (
	.clk(clk),
	.d(\WideOr7~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_0),
	.prn(vcc));
defparam \master_address[0] .is_wysiwyg = "true";
defparam \master_address[0] .power_up = "low";

dffeas \master_address[1] (
	.clk(clk),
	.d(\WideOr6~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_1),
	.prn(vcc));
defparam \master_address[1] .is_wysiwyg = "true";
defparam \master_address[1] .power_up = "low";

dffeas master_read(
	.clk(clk),
	.d(\WideOr9~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_read1),
	.prn(vcc));
defparam master_read.is_wysiwyg = "true";
defparam master_read.power_up = "low";

dffeas \readdata_for_user[2] (
	.clk(clk),
	.d(basic_reconfig_readdata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_2),
	.prn(vcc));
defparam \readdata_for_user[2] .is_wysiwyg = "true";
defparam \readdata_for_user[2] .power_up = "low";

dffeas \readdata_for_user[0] (
	.clk(clk),
	.d(basic_reconfig_readdata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_0),
	.prn(vcc));
defparam \readdata_for_user[0] .is_wysiwyg = "true";
defparam \readdata_for_user[0] .power_up = "low";

dffeas \readdata_for_user[3] (
	.clk(clk),
	.d(basic_reconfig_readdata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_3),
	.prn(vcc));
defparam \readdata_for_user[3] .is_wysiwyg = "true";
defparam \readdata_for_user[3] .power_up = "low";

dffeas \readdata_for_user[1] (
	.clk(clk),
	.d(basic_reconfig_readdata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_1),
	.prn(vcc));
defparam \readdata_for_user[1] .is_wysiwyg = "true";
defparam \readdata_for_user[1] .power_up = "low";

dffeas \readdata_for_user[10] (
	.clk(clk),
	.d(basic_reconfig_readdata_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_10),
	.prn(vcc));
defparam \readdata_for_user[10] .is_wysiwyg = "true";
defparam \readdata_for_user[10] .power_up = "low";

dffeas \readdata_for_user[8] (
	.clk(clk),
	.d(basic_reconfig_readdata_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_8),
	.prn(vcc));
defparam \readdata_for_user[8] .is_wysiwyg = "true";
defparam \readdata_for_user[8] .power_up = "low";

dffeas \readdata_for_user[11] (
	.clk(clk),
	.d(basic_reconfig_readdata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_11),
	.prn(vcc));
defparam \readdata_for_user[11] .is_wysiwyg = "true";
defparam \readdata_for_user[11] .power_up = "low";

dffeas \readdata_for_user[9] (
	.clk(clk),
	.d(basic_reconfig_readdata_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_9),
	.prn(vcc));
defparam \readdata_for_user[9] .is_wysiwyg = "true";
defparam \readdata_for_user[9] .power_up = "low";

dffeas \readdata_for_user[6] (
	.clk(clk),
	.d(basic_reconfig_readdata_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_6),
	.prn(vcc));
defparam \readdata_for_user[6] .is_wysiwyg = "true";
defparam \readdata_for_user[6] .power_up = "low";

dffeas \readdata_for_user[4] (
	.clk(clk),
	.d(basic_reconfig_readdata_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_4),
	.prn(vcc));
defparam \readdata_for_user[4] .is_wysiwyg = "true";
defparam \readdata_for_user[4] .power_up = "low";

dffeas \readdata_for_user[7] (
	.clk(clk),
	.d(basic_reconfig_readdata_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_7),
	.prn(vcc));
defparam \readdata_for_user[7] .is_wysiwyg = "true";
defparam \readdata_for_user[7] .power_up = "low";

dffeas \readdata_for_user[5] (
	.clk(clk),
	.d(basic_reconfig_readdata_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_5),
	.prn(vcc));
defparam \readdata_for_user[5] .is_wysiwyg = "true";
defparam \readdata_for_user[5] .power_up = "low";

dffeas \readdata_for_user[14] (
	.clk(clk),
	.d(basic_reconfig_readdata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_14),
	.prn(vcc));
defparam \readdata_for_user[14] .is_wysiwyg = "true";
defparam \readdata_for_user[14] .power_up = "low";

dffeas \readdata_for_user[12] (
	.clk(clk),
	.d(basic_reconfig_readdata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_12),
	.prn(vcc));
defparam \readdata_for_user[12] .is_wysiwyg = "true";
defparam \readdata_for_user[12] .power_up = "low";

dffeas \readdata_for_user[15] (
	.clk(clk),
	.d(basic_reconfig_readdata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_15),
	.prn(vcc));
defparam \readdata_for_user[15] .is_wysiwyg = "true";
defparam \readdata_for_user[15] .power_up = "low";

dffeas \readdata_for_user[13] (
	.clk(clk),
	.d(basic_reconfig_readdata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_13),
	.prn(vcc));
defparam \readdata_for_user[13] .is_wysiwyg = "true";
defparam \readdata_for_user[13] .power_up = "low";

dffeas \readdata_for_user[16] (
	.clk(clk),
	.d(basic_reconfig_readdata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_16),
	.prn(vcc));
defparam \readdata_for_user[16] .is_wysiwyg = "true";
defparam \readdata_for_user[16] .power_up = "low";

dffeas \ph_readdata[0] (
	.clk(clk),
	.d(basic_reconfig_readdata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_0),
	.prn(vcc));
defparam \ph_readdata[0] .is_wysiwyg = "true";
defparam \ph_readdata[0] .power_up = "low";

dffeas \ph_readdata[1] (
	.clk(clk),
	.d(basic_reconfig_readdata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_1),
	.prn(vcc));
defparam \ph_readdata[1] .is_wysiwyg = "true";
defparam \ph_readdata[1] .power_up = "low";

dffeas \readdata_for_user[17] (
	.clk(clk),
	.d(basic_reconfig_readdata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_17),
	.prn(vcc));
defparam \readdata_for_user[17] .is_wysiwyg = "true";
defparam \readdata_for_user[17] .power_up = "low";

dffeas \ph_readdata[2] (
	.clk(clk),
	.d(basic_reconfig_readdata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_2),
	.prn(vcc));
defparam \ph_readdata[2] .is_wysiwyg = "true";
defparam \ph_readdata[2] .power_up = "low";

dffeas \readdata_for_user[18] (
	.clk(clk),
	.d(basic_reconfig_readdata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_18),
	.prn(vcc));
defparam \readdata_for_user[18] .is_wysiwyg = "true";
defparam \readdata_for_user[18] .power_up = "low";

dffeas \ph_readdata[3] (
	.clk(clk),
	.d(basic_reconfig_readdata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_3),
	.prn(vcc));
defparam \ph_readdata[3] .is_wysiwyg = "true";
defparam \ph_readdata[3] .power_up = "low";

dffeas \readdata_for_user[19] (
	.clk(clk),
	.d(basic_reconfig_readdata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_19),
	.prn(vcc));
defparam \readdata_for_user[19] .is_wysiwyg = "true";
defparam \readdata_for_user[19] .power_up = "low";

dffeas \ph_readdata[4] (
	.clk(clk),
	.d(basic_reconfig_readdata_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_4),
	.prn(vcc));
defparam \ph_readdata[4] .is_wysiwyg = "true";
defparam \ph_readdata[4] .power_up = "low";

dffeas \readdata_for_user[20] (
	.clk(clk),
	.d(basic_reconfig_readdata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_20),
	.prn(vcc));
defparam \readdata_for_user[20] .is_wysiwyg = "true";
defparam \readdata_for_user[20] .power_up = "low";

dffeas \ph_readdata[5] (
	.clk(clk),
	.d(basic_reconfig_readdata_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_5),
	.prn(vcc));
defparam \ph_readdata[5] .is_wysiwyg = "true";
defparam \ph_readdata[5] .power_up = "low";

dffeas \readdata_for_user[21] (
	.clk(clk),
	.d(basic_reconfig_readdata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_21),
	.prn(vcc));
defparam \readdata_for_user[21] .is_wysiwyg = "true";
defparam \readdata_for_user[21] .power_up = "low";

dffeas \ph_readdata[6] (
	.clk(clk),
	.d(basic_reconfig_readdata_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_6),
	.prn(vcc));
defparam \ph_readdata[6] .is_wysiwyg = "true";
defparam \ph_readdata[6] .power_up = "low";

dffeas \readdata_for_user[22] (
	.clk(clk),
	.d(basic_reconfig_readdata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_22),
	.prn(vcc));
defparam \readdata_for_user[22] .is_wysiwyg = "true";
defparam \readdata_for_user[22] .power_up = "low";

dffeas \ph_readdata[7] (
	.clk(clk),
	.d(basic_reconfig_readdata_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_7),
	.prn(vcc));
defparam \ph_readdata[7] .is_wysiwyg = "true";
defparam \ph_readdata[7] .power_up = "low";

dffeas \readdata_for_user[23] (
	.clk(clk),
	.d(basic_reconfig_readdata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_23),
	.prn(vcc));
defparam \readdata_for_user[23] .is_wysiwyg = "true";
defparam \readdata_for_user[23] .power_up = "low";

dffeas \ph_readdata[8] (
	.clk(clk),
	.d(basic_reconfig_readdata_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_8),
	.prn(vcc));
defparam \ph_readdata[8] .is_wysiwyg = "true";
defparam \ph_readdata[8] .power_up = "low";

dffeas \readdata_for_user[24] (
	.clk(clk),
	.d(basic_reconfig_readdata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_24),
	.prn(vcc));
defparam \readdata_for_user[24] .is_wysiwyg = "true";
defparam \readdata_for_user[24] .power_up = "low";

dffeas \ph_readdata[9] (
	.clk(clk),
	.d(basic_reconfig_readdata_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_9),
	.prn(vcc));
defparam \ph_readdata[9] .is_wysiwyg = "true";
defparam \ph_readdata[9] .power_up = "low";

dffeas \ph_readdata[10] (
	.clk(clk),
	.d(basic_reconfig_readdata_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_10),
	.prn(vcc));
defparam \ph_readdata[10] .is_wysiwyg = "true";
defparam \ph_readdata[10] .power_up = "low";

dffeas \readdata_for_user[25] (
	.clk(clk),
	.d(basic_reconfig_readdata_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_25),
	.prn(vcc));
defparam \readdata_for_user[25] .is_wysiwyg = "true";
defparam \readdata_for_user[25] .power_up = "low";

dffeas \ph_readdata[11] (
	.clk(clk),
	.d(basic_reconfig_readdata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_11),
	.prn(vcc));
defparam \ph_readdata[11] .is_wysiwyg = "true";
defparam \ph_readdata[11] .power_up = "low";

dffeas \readdata_for_user[26] (
	.clk(clk),
	.d(basic_reconfig_readdata_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_26),
	.prn(vcc));
defparam \readdata_for_user[26] .is_wysiwyg = "true";
defparam \readdata_for_user[26] .power_up = "low";

dffeas \ph_readdata[12] (
	.clk(clk),
	.d(basic_reconfig_readdata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_12),
	.prn(vcc));
defparam \ph_readdata[12] .is_wysiwyg = "true";
defparam \ph_readdata[12] .power_up = "low";

dffeas \readdata_for_user[27] (
	.clk(clk),
	.d(basic_reconfig_readdata_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_27),
	.prn(vcc));
defparam \readdata_for_user[27] .is_wysiwyg = "true";
defparam \readdata_for_user[27] .power_up = "low";

dffeas \ph_readdata[13] (
	.clk(clk),
	.d(basic_reconfig_readdata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_13),
	.prn(vcc));
defparam \ph_readdata[13] .is_wysiwyg = "true";
defparam \ph_readdata[13] .power_up = "low";

dffeas \readdata_for_user[28] (
	.clk(clk),
	.d(basic_reconfig_readdata_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_28),
	.prn(vcc));
defparam \readdata_for_user[28] .is_wysiwyg = "true";
defparam \readdata_for_user[28] .power_up = "low";

dffeas \ph_readdata[14] (
	.clk(clk),
	.d(basic_reconfig_readdata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_14),
	.prn(vcc));
defparam \ph_readdata[14] .is_wysiwyg = "true";
defparam \ph_readdata[14] .power_up = "low";

dffeas \readdata_for_user[29] (
	.clk(clk),
	.d(basic_reconfig_readdata_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_29),
	.prn(vcc));
defparam \readdata_for_user[29] .is_wysiwyg = "true";
defparam \readdata_for_user[29] .power_up = "low";

dffeas \ph_readdata[15] (
	.clk(clk),
	.d(basic_reconfig_readdata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_15),
	.prn(vcc));
defparam \ph_readdata[15] .is_wysiwyg = "true";
defparam \ph_readdata[15] .power_up = "low";

dffeas \readdata_for_user[30] (
	.clk(clk),
	.d(basic_reconfig_readdata_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_30),
	.prn(vcc));
defparam \readdata_for_user[30] .is_wysiwyg = "true";
defparam \readdata_for_user[30] .power_up = "low";

dffeas \ph_readdata[16] (
	.clk(clk),
	.d(basic_reconfig_readdata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_16),
	.prn(vcc));
defparam \ph_readdata[16] .is_wysiwyg = "true";
defparam \ph_readdata[16] .power_up = "low";

dffeas \readdata_for_user[31] (
	.clk(clk),
	.d(basic_reconfig_readdata_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_31),
	.prn(vcc));
defparam \readdata_for_user[31] .is_wysiwyg = "true";
defparam \readdata_for_user[31] .power_up = "low";

dffeas \ph_readdata[17] (
	.clk(clk),
	.d(basic_reconfig_readdata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_17),
	.prn(vcc));
defparam \ph_readdata[17] .is_wysiwyg = "true";
defparam \ph_readdata[17] .power_up = "low";

dffeas \ph_readdata[18] (
	.clk(clk),
	.d(basic_reconfig_readdata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_18),
	.prn(vcc));
defparam \ph_readdata[18] .is_wysiwyg = "true";
defparam \ph_readdata[18] .power_up = "low";

dffeas \ph_readdata[19] (
	.clk(clk),
	.d(basic_reconfig_readdata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_19),
	.prn(vcc));
defparam \ph_readdata[19] .is_wysiwyg = "true";
defparam \ph_readdata[19] .power_up = "low";

dffeas \ph_readdata[20] (
	.clk(clk),
	.d(basic_reconfig_readdata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_20),
	.prn(vcc));
defparam \ph_readdata[20] .is_wysiwyg = "true";
defparam \ph_readdata[20] .power_up = "low";

dffeas \ph_readdata[21] (
	.clk(clk),
	.d(basic_reconfig_readdata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_21),
	.prn(vcc));
defparam \ph_readdata[21] .is_wysiwyg = "true";
defparam \ph_readdata[21] .power_up = "low";

dffeas \ph_readdata[22] (
	.clk(clk),
	.d(basic_reconfig_readdata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_22),
	.prn(vcc));
defparam \ph_readdata[22] .is_wysiwyg = "true";
defparam \ph_readdata[22] .power_up = "low";

dffeas \ph_readdata[23] (
	.clk(clk),
	.d(basic_reconfig_readdata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_23),
	.prn(vcc));
defparam \ph_readdata[23] .is_wysiwyg = "true";
defparam \ph_readdata[23] .power_up = "low";

dffeas \ph_readdata[24] (
	.clk(clk),
	.d(basic_reconfig_readdata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_24),
	.prn(vcc));
defparam \ph_readdata[24] .is_wysiwyg = "true";
defparam \ph_readdata[24] .power_up = "low";

dffeas \ph_readdata[25] (
	.clk(clk),
	.d(basic_reconfig_readdata_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_25),
	.prn(vcc));
defparam \ph_readdata[25] .is_wysiwyg = "true";
defparam \ph_readdata[25] .power_up = "low";

dffeas \ph_readdata[26] (
	.clk(clk),
	.d(basic_reconfig_readdata_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_26),
	.prn(vcc));
defparam \ph_readdata[26] .is_wysiwyg = "true";
defparam \ph_readdata[26] .power_up = "low";

dffeas \ph_readdata[27] (
	.clk(clk),
	.d(basic_reconfig_readdata_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_27),
	.prn(vcc));
defparam \ph_readdata[27] .is_wysiwyg = "true";
defparam \ph_readdata[27] .power_up = "low";

dffeas \ph_readdata[28] (
	.clk(clk),
	.d(basic_reconfig_readdata_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_28),
	.prn(vcc));
defparam \ph_readdata[28] .is_wysiwyg = "true";
defparam \ph_readdata[28] .power_up = "low";

dffeas \ph_readdata[29] (
	.clk(clk),
	.d(basic_reconfig_readdata_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_29),
	.prn(vcc));
defparam \ph_readdata[29] .is_wysiwyg = "true";
defparam \ph_readdata[29] .power_up = "low";

dffeas \ph_readdata[30] (
	.clk(clk),
	.d(basic_reconfig_readdata_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_30),
	.prn(vcc));
defparam \ph_readdata[30] .is_wysiwyg = "true";
defparam \ph_readdata[30] .power_up = "low";

dffeas \ph_readdata[31] (
	.clk(clk),
	.d(basic_reconfig_readdata_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(ph_readdata_31),
	.prn(vcc));
defparam \ph_readdata[31] .is_wysiwyg = "true";
defparam \ph_readdata[31] .power_up = "low";

dffeas \master_writedata[1] (
	.clk(clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_1),
	.prn(vcc));
defparam \master_writedata[1] .is_wysiwyg = "true";
defparam \master_writedata[1] .power_up = "low";

dffeas \master_writedata[2] (
	.clk(clk),
	.d(\Selector25~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_2),
	.prn(vcc));
defparam \master_writedata[2] .is_wysiwyg = "true";
defparam \master_writedata[2] .power_up = "low";

dffeas \master_writedata[0] (
	.clk(clk),
	.d(\Selector27~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_0),
	.prn(vcc));
defparam \master_writedata[0] .is_wysiwyg = "true";
defparam \master_writedata[0] .power_up = "low";

dffeas \master_writedata[3] (
	.clk(clk),
	.d(\Selector24~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_3),
	.prn(vcc));
defparam \master_writedata[3] .is_wysiwyg = "true";
defparam \master_writedata[3] .power_up = "low";

dffeas \master_writedata[4] (
	.clk(clk),
	.d(\Selector23~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_4),
	.prn(vcc));
defparam \master_writedata[4] .is_wysiwyg = "true";
defparam \master_writedata[4] .power_up = "low";

dffeas \master_writedata[5] (
	.clk(clk),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_5),
	.prn(vcc));
defparam \master_writedata[5] .is_wysiwyg = "true";
defparam \master_writedata[5] .power_up = "low";

dffeas \master_writedata[6] (
	.clk(clk),
	.d(\Selector21~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_6),
	.prn(vcc));
defparam \master_writedata[6] .is_wysiwyg = "true";
defparam \master_writedata[6] .power_up = "low";

dffeas \master_writedata[7] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_7),
	.prn(vcc));
defparam \master_writedata[7] .is_wysiwyg = "true";
defparam \master_writedata[7] .power_up = "low";

dffeas \master_writedata[8] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_8),
	.prn(vcc));
defparam \master_writedata[8] .is_wysiwyg = "true";
defparam \master_writedata[8] .power_up = "low";

dffeas \master_writedata[9] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_9),
	.prn(vcc));
defparam \master_writedata[9] .is_wysiwyg = "true";
defparam \master_writedata[9] .power_up = "low";

dffeas \master_writedata[10] (
	.clk(clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_10),
	.prn(vcc));
defparam \master_writedata[10] .is_wysiwyg = "true";
defparam \master_writedata[10] .power_up = "low";

dffeas waitrequest_to_ctrl(
	.clk(clk),
	.d(\Selector16~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_to_ctrl1),
	.prn(vcc));
defparam waitrequest_to_ctrl.is_wysiwyg = "true";
defparam waitrequest_to_ctrl.power_up = "low";

dffeas illegal_phy_ch(
	.clk(clk),
	.d(Equal8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[6]~0_combout ),
	.q(illegal_phy_ch1),
	.prn(vcc));
defparam illegal_phy_ch.is_wysiwyg = "true";
defparam illegal_phy_ch.power_up = "low";

dffeas \lch_dly[7] (
	.clk(clk),
	.d(logical_ch_addr[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[7]~q ),
	.prn(vcc));
defparam \lch_dly[7] .is_wysiwyg = "true";
defparam \lch_dly[7] .power_up = "low";

dffeas \lch_dly[5] (
	.clk(clk),
	.d(logical_ch_addr[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[5]~q ),
	.prn(vcc));
defparam \lch_dly[5] .is_wysiwyg = "true";
defparam \lch_dly[5] .power_up = "low";

dffeas \lch_dly[6] (
	.clk(clk),
	.d(logical_ch_addr[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[6]~q ),
	.prn(vcc));
defparam \lch_dly[6] .is_wysiwyg = "true";
defparam \lch_dly[6] .power_up = "low";

cyclonev_lcell_comb \lch_legal~0 (
	.dataa(!logical_ch_addr[5]),
	.datab(!logical_ch_addr[6]),
	.datac(!\lch_dly[5]~q ),
	.datad(!\lch_dly[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~0 .extended_lut = "off";
defparam \lch_legal~0 .lut_mask = 64'h8421842184218421;
defparam \lch_legal~0 .shared_arith = "off";

dffeas \lch_dly[8] (
	.clk(clk),
	.d(logical_ch_addr[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[8]~q ),
	.prn(vcc));
defparam \lch_dly[8] .is_wysiwyg = "true";
defparam \lch_dly[8] .power_up = "low";

dffeas \lch_dly[9] (
	.clk(clk),
	.d(logical_ch_addr[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[9]~q ),
	.prn(vcc));
defparam \lch_dly[9] .is_wysiwyg = "true";
defparam \lch_dly[9] .power_up = "low";

cyclonev_lcell_comb \lch_legal~1 (
	.dataa(!logical_ch_addr[8]),
	.datab(!logical_ch_addr[9]),
	.datac(!\lch_dly[8]~q ),
	.datad(!\lch_dly[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~1 .extended_lut = "off";
defparam \lch_legal~1 .lut_mask = 64'h8421842184218421;
defparam \lch_legal~1 .shared_arith = "off";

dffeas \lch_dly[4] (
	.clk(clk),
	.d(logical_ch_addr[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[4]~q ),
	.prn(vcc));
defparam \lch_dly[4] .is_wysiwyg = "true";
defparam \lch_dly[4] .power_up = "low";

cyclonev_lcell_comb \Selector5~2 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~2 .extended_lut = "off";
defparam \Selector5~2 .lut_mask = 64'h4444444444444444;
defparam \Selector5~2 .shared_arith = "off";

dffeas \lch_dly[0] (
	.clk(clk),
	.d(logical_ch_addr[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[0]~q ),
	.prn(vcc));
defparam \lch_dly[0] .is_wysiwyg = "true";
defparam \lch_dly[0] .power_up = "low";

dffeas \lch_dly[1] (
	.clk(clk),
	.d(logical_ch_addr[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[1]~q ),
	.prn(vcc));
defparam \lch_dly[1] .is_wysiwyg = "true";
defparam \lch_dly[1] .power_up = "low";

cyclonev_lcell_comb \lch_legal~2 (
	.dataa(!logical_ch_addr[0]),
	.datab(!logical_ch_addr[1]),
	.datac(!\Selector5~2_combout ),
	.datad(!\lch_dly[0]~q ),
	.datae(!\lch_dly[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~2 .extended_lut = "off";
defparam \lch_legal~2 .lut_mask = 64'h8040201080402010;
defparam \lch_legal~2 .shared_arith = "off";

dffeas \lch_dly[2] (
	.clk(clk),
	.d(logical_ch_addr[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[2]~q ),
	.prn(vcc));
defparam \lch_dly[2] .is_wysiwyg = "true";
defparam \lch_dly[2] .power_up = "low";

dffeas \lch_dly[3] (
	.clk(clk),
	.d(logical_ch_addr[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[3]~q ),
	.prn(vcc));
defparam \lch_dly[3] .is_wysiwyg = "true";
defparam \lch_dly[3] .power_up = "low";

cyclonev_lcell_comb \lch_legal~3 (
	.dataa(!logical_ch_addr[2]),
	.datab(!logical_ch_addr[3]),
	.datac(!\lch_dly[2]~q ),
	.datad(!\lch_dly[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~3 .extended_lut = "off";
defparam \lch_legal~3 .lut_mask = 64'h8421842184218421;
defparam \lch_legal~3 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~4 (
	.dataa(!logical_ch_addr[4]),
	.datab(!\lch_dly[4]~q ),
	.datac(!\lch_legal~2_combout ),
	.datad(!\lch_legal~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~4 .extended_lut = "off";
defparam \lch_legal~4 .lut_mask = 64'h0009000900090009;
defparam \lch_legal~4 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~5 (
	.dataa(!logical_ch_addr[7]),
	.datab(!\lch_dly[7]~q ),
	.datac(!\lch_legal~0_combout ),
	.datad(!\lch_legal~1_combout ),
	.datae(!\lch_legal~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~5 .extended_lut = "off";
defparam \lch_legal~5 .lut_mask = 64'h0000000900000009;
defparam \lch_legal~5 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~6 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!Equal8),
	.datad(!\lch_legal~q ),
	.datae(!\lch_legal~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~6 .extended_lut = "off";
defparam \lch_legal~6 .lut_mask = 64'h000020FF000020FF;
defparam \lch_legal~6 .shared_arith = "off";

dffeas lch_legal(
	.clk(clk),
	.d(\lch_legal~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_legal~q ),
	.prn(vcc));
defparam lch_legal.is_wysiwyg = "true";
defparam lch_legal.power_up = "low";

dffeas \state.ST_WRITE_DATA_TO_RECONFIG_BASIC (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.prn(vcc));
defparam \state.ST_WRITE_DATA_TO_RECONFIG_BASIC .is_wysiwyg = "true";
defparam \state.ST_WRITE_DATA_TO_RECONFIG_BASIC .power_up = "low";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.dataf(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h00007FFF8000FFFF;
defparam \Selector9~0 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_WRITE (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_WRITE .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_WRITE .power_up = "low";

cyclonev_lcell_comb \Selector6~1 (
	.dataa(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datab(!Equal8),
	.datac(!\lch_legal~q ),
	.datad(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datae(!\Selector5~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'h444F000F444F000F;
defparam \Selector6~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~2 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.datae(!\Selector6~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~2 .extended_lut = "off";
defparam \Selector6~2 .lut_mask = 64'h00FB0CFF00FB0CFF;
defparam \Selector6~2 .shared_arith = "off";

dffeas \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK (
	.clk(clk),
	.d(\Selector6~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.prn(vcc));
defparam \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK .is_wysiwyg = "true";
defparam \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK .power_up = "low";

cyclonev_lcell_comb \Selector13~0 (
	.dataa(!ctrl_go),
	.datab(!\state.ST_START_AGAIN~q ),
	.datac(!ctrl_lock),
	.datad(!\state.ST_CHECK_CTRLLOCK~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~0 .extended_lut = "off";
defparam \Selector13~0 .lut_mask = 64'h222F222F222F222F;
defparam \Selector13~0 .shared_arith = "off";

dffeas \state.ST_START_AGAIN (
	.clk(clk),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_START_AGAIN~q ),
	.prn(vcc));
defparam \state.ST_START_AGAIN .is_wysiwyg = "true";
defparam \state.ST_START_AGAIN .power_up = "low";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!ctrl_go),
	.datab(!\state.ST_START_AGAIN~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h1111111111111111;
defparam \Selector7~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~1 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!basic_reconfig_waitrequest2),
	.datac(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datad(!\Selector5~2_combout ),
	.datae(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.dataf(!\Selector7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~1 .extended_lut = "off";
defparam \Selector7~1 .lut_mask = 64'h030F474FFFFFFFFF;
defparam \Selector7~1 .shared_arith = "off";

dffeas \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG (
	.clk(clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.prn(vcc));
defparam \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG .is_wysiwyg = "true";
defparam \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG .power_up = "low";

cyclonev_lcell_comb \Selector5~4 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.dataf(!\Selector5~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~4 .extended_lut = "off";
defparam \Selector5~4 .lut_mask = 64'h0000800000000000;
defparam \Selector5~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~5 (
	.dataa(!\lch_legal~q ),
	.datab(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datac(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~5 .extended_lut = "off";
defparam \Selector5~5 .lut_mask = 64'h0D0D0D0D0D0D0D0D;
defparam \Selector5~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~6 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector5~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~6 .extended_lut = "off";
defparam \Selector5~6 .lut_mask = 64'h8000000080000000;
defparam \Selector5~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~7 (
	.dataa(!\state.0000~q ),
	.datab(!\state.ST_REQ_MUTEX~q ),
	.datac(!\state.ST_START_AGAIN~q ),
	.datad(!\state.ST_CHECK_CTRLLOCK~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~7 .extended_lut = "off";
defparam \Selector5~7 .lut_mask = 64'h4000400040004000;
defparam \Selector5~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!\Selector5~3_combout ),
	.datab(!ctrl_opcode_0),
	.datac(!\Selector5~4_combout ),
	.datad(!\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.datae(!\Selector5~6_combout ),
	.dataf(!\Selector5~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h0C0C0C0C0CAC0C0C;
defparam \Selector10~0 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_READ (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_READ .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_READ .power_up = "low";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.dataf(!\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h00007FFF8000FFFF;
defparam \Selector11~0 .shared_arith = "off";

dffeas \state.ST_READ_RECONFIG_BASIC_DATA (
	.clk(clk),
	.d(\Selector11~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.prn(vcc));
defparam \state.ST_READ_RECONFIG_BASIC_DATA .is_wysiwyg = "true";
defparam \state.ST_READ_RECONFIG_BASIC_DATA .power_up = "low";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.datab(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'h8888888888888888;
defparam \Selector12~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~1 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!Equal8),
	.datad(!\state.ST_CHECK_CTRLLOCK~q ),
	.datae(!\Selector5~2_combout ),
	.dataf(!\Selector12~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~1 .extended_lut = "off";
defparam \Selector12~1 .lut_mask = 64'hAAFFAAFF00002020;
defparam \Selector12~1 .shared_arith = "off";

dffeas \state.ST_CHECK_CTRLLOCK (
	.clk(clk),
	.d(\Selector12~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CHECK_CTRLLOCK~q ),
	.prn(vcc));
defparam \state.ST_CHECK_CTRLLOCK .is_wysiwyg = "true";
defparam \state.ST_CHECK_CTRLLOCK .power_up = "low";

cyclonev_lcell_comb \Selector14~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_RELEASE_REQ~q ),
	.datad(!ctrl_lock),
	.datae(!\state.ST_CHECK_CTRLLOCK~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~0 .extended_lut = "off";
defparam \Selector14~0 .lut_mask = 64'h0D0DFF0D0D0DFF0D;
defparam \Selector14~0 .shared_arith = "off";

dffeas \state.ST_RELEASE_REQ (
	.clk(clk),
	.d(\Selector14~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_RELEASE_REQ~q ),
	.prn(vcc));
defparam \state.ST_RELEASE_REQ .is_wysiwyg = "true";
defparam \state.ST_RELEASE_REQ .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_RELEASE_REQ~q ),
	.datad(!\Selector5~3_combout ),
	.datae(!ctrl_go),
	.dataf(!\state.0000~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h0000FD00FD00FD00;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.0000 (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.0000~q ),
	.prn(vcc));
defparam \state.0000 .is_wysiwyg = "true";
defparam \state.0000 .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!mutex_grant),
	.datab(!ctrl_go),
	.datac(!\state.0000~q ),
	.datad(!\state.ST_REQ_MUTEX~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h30BA30BA30BA30BA;
defparam \Selector1~0 .shared_arith = "off";

dffeas \state.ST_REQ_MUTEX (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_REQ_MUTEX~q ),
	.prn(vcc));
defparam \state.ST_REQ_MUTEX .is_wysiwyg = "true";
defparam \state.ST_REQ_MUTEX .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!mutex_grant),
	.datab(!\state.ST_REQ_MUTEX~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h1111111111111111;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h00007FFFFFFFFFFF;
defparam \Selector2~1 .shared_arith = "off";

dffeas \state.ST_WRITE_RECONFIG_BASIC_LCH (
	.clk(clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.prn(vcc));
defparam \state.ST_WRITE_RECONFIG_BASIC_LCH .is_wysiwyg = "true";
defparam \state.ST_WRITE_RECONFIG_BASIC_LCH .power_up = "low";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\Selector5~3_combout ),
	.datac(!\state.ST_READ_PHY_ADDRESS~q ),
	.datad(!\lch_legal~q ),
	.datae(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.dataf(!\Selector5~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h04048C0400000000;
defparam \Selector3~0 .shared_arith = "off";

dffeas \state.ST_READ_PHY_ADDRESS (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_READ_PHY_ADDRESS~q ),
	.prn(vcc));
defparam \state.ST_READ_PHY_ADDRESS .is_wysiwyg = "true";
defparam \state.ST_READ_PHY_ADDRESS .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!Equal8),
	.datad(!\state.ST_READ_PHY_ADDRESS~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h10BA10BA10BA10BA;
defparam \Selector4~0 .shared_arith = "off";

dffeas \state.ST_CHECK_PHY_ADD_LEGAL (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.prn(vcc));
defparam \state.ST_CHECK_PHY_ADD_LEGAL .is_wysiwyg = "true";
defparam \state.ST_CHECK_PHY_ADD_LEGAL .power_up = "low";

cyclonev_lcell_comb \Selector5~3 (
	.dataa(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datab(!Equal8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~3 .extended_lut = "off";
defparam \Selector5~3 .lut_mask = 64'h1111111111111111;
defparam \Selector5~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!\Selector5~3_combout ),
	.datab(!ctrl_opcode_0),
	.datac(!\Selector5~4_combout ),
	.datad(!\Selector5~6_combout ),
	.datae(!\Selector5~7_combout ),
	.dataf(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h030303030303A303;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr7~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\Selector13~0_combout ),
	.datac(!\Selector3~0_combout ),
	.datad(!\Selector4~0_combout ),
	.datae(!\Selector12~1_combout ),
	.dataf(!\Selector0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr7~0 .extended_lut = "off";
defparam \WideOr7~0 .lut_mask = 64'h0000000080000000;
defparam \WideOr7~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr8(
	.dataa(!\Selector11~0_combout ),
	.datab(!\Selector6~2_combout ),
	.datac(!\WideOr7~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr8~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr8.extended_lut = "off";
defparam WideOr8.lut_mask = 64'h0808080808080808;
defparam WideOr8.shared_arith = "off";

cyclonev_lcell_comb \WideOr5~0 (
	.dataa(!\Selector11~0_combout ),
	.datab(!\Selector8~0_combout ),
	.datac(!\Selector7~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr5~0 .extended_lut = "off";
defparam \WideOr5~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \WideOr5~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr17~0 (
	.dataa(!\Selector13~0_combout ),
	.datab(!\Selector3~0_combout ),
	.datac(!\Selector6~2_combout ),
	.datad(!\Selector2~1_combout ),
	.datae(!\Selector10~0_combout ),
	.dataf(!\Selector9~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~0 .extended_lut = "off";
defparam \WideOr17~0 .lut_mask = 64'h8000000000000000;
defparam \WideOr17~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!mutex_req1),
	.datab(!\Selector1~0_combout ),
	.datac(!\Selector4~0_combout ),
	.datad(!\Selector12~1_combout ),
	.datae(!\WideOr5~0_combout ),
	.dataf(!\WideOr17~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h7777777737777777;
defparam \Selector28~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr7(
	.dataa(!\WideOr7~0_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr7~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr7.extended_lut = "off";
defparam WideOr7.lut_mask = 64'h4444444444444444;
defparam WideOr7.shared_arith = "off";

cyclonev_lcell_comb WideOr6(
	.dataa(!\Selector3~0_combout ),
	.datab(!\Selector6~2_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Selector9~0_combout ),
	.datae(!\Selector14~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr6~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr6.extended_lut = "off";
defparam WideOr6.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr6.shared_arith = "off";

cyclonev_lcell_comb WideOr9(
	.dataa(!\Selector3~0_combout ),
	.datab(!\Selector11~0_combout ),
	.datac(!\Selector6~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr9~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr9.extended_lut = "off";
defparam WideOr9.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam WideOr9.shared_arith = "off";

cyclonev_lcell_comb \Selector12~2 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datad(!Equal8),
	.datae(!\Selector5~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~2 .extended_lut = "off";
defparam \Selector12~2 .lut_mask = 64'h0000020000000200;
defparam \Selector12~2 .shared_arith = "off";

cyclonev_lcell_comb \readdata_for_user[0]~0 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\state.ST_CHECK_CTRLLOCK~q ),
	.datac(!\Selector12~2_combout ),
	.datad(gnd),
	.datae(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata_for_user[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata_for_user[0]~0 .extended_lut = "off";
defparam \readdata_for_user[0]~0 .lut_mask = 64'h0000BFBF0000BFBF;
defparam \readdata_for_user[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_RELEASE_REQ~q ),
	.datad(!\Selector1~0_combout ),
	.datae(!ctrl_lock),
	.dataf(!\state.ST_CHECK_CTRLLOCK~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'hF200F2000000F200;
defparam \Selector16~0 .shared_arith = "off";

cyclonev_lcell_comb \ph_readdata[6]~0 (
	.dataa(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datab(!\Selector12~1_combout ),
	.datac(!\Selector0~0_combout ),
	.datad(!\WideOr5~0_combout ),
	.datae(!\WideOr17~0_combout ),
	.dataf(!\Selector16~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ph_readdata[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ph_readdata[6]~0 .extended_lut = "off";
defparam \ph_readdata[6]~0 .lut_mask = 64'h0000000000000D00;
defparam \ph_readdata[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!uif_addr_offset_1),
	.datae(!Decoder3),
	.dataf(!lpbk_lock),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'h0000628000006680;
defparam \Selector26~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~1 (
	.dataa(!logical_ch_addr[1]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!\Selector7~1_combout ),
	.datae(!outdata_1),
	.dataf(!\Selector26~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~1 .extended_lut = "off";
defparam \Selector26~1 .lut_mask = 64'h11111F1F11FF1FFF;
defparam \Selector26~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!logical_ch_addr[2]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector14~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \Selector25~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~1 (
	.dataa(!uif_addr_offset_1),
	.datab(!analog_length),
	.datac(!\Selector8~0_combout ),
	.datad(!\Selector7~1_combout ),
	.datae(!outdata_2),
	.dataf(!\Selector25~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~1 .extended_lut = "off";
defparam \Selector25~1 .lut_mask = 64'hFFFFFFFF00220F2F;
defparam \Selector25~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_0),
	.datad(!uif_addr_offset_1),
	.datae(!Decoder3),
	.dataf(!lpbk_lock),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h0000628000002080;
defparam \Selector27~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~1 (
	.dataa(!logical_ch_addr[0]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~1 .extended_lut = "off";
defparam \Selector27~1 .lut_mask = 64'h111F111F111F111F;
defparam \Selector27~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~2 (
	.dataa(!\Selector10~0_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(!\Selector27~0_combout ),
	.datad(!\Selector27~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~2 .extended_lut = "off";
defparam \Selector27~2 .lut_mask = 64'h57FF57FF57FF57FF;
defparam \Selector27~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_0),
	.datac(!\Selector9~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h0101010101010101;
defparam \Selector24~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~1 (
	.dataa(!logical_ch_addr[3]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_3),
	.datae(!\Selector24~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~1 .extended_lut = "off";
defparam \Selector24~1 .lut_mask = 64'h111FFFFF111FFFFF;
defparam \Selector24~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector23~0 (
	.dataa(!logical_ch_addr[4]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h111F111F111F111F;
defparam \Selector23~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector23~1 (
	.dataa(!uif_addr_offset_3),
	.datab(!\Selector7~1_combout ),
	.datac(!WideOr5),
	.datad(!\Selector23~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~1 .extended_lut = "off";
defparam \Selector23~1 .lut_mask = 64'h02FF02FF02FF02FF;
defparam \Selector23~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector22~0 (
	.dataa(!logical_ch_addr[5]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector22~0 .extended_lut = "off";
defparam \Selector22~0 .lut_mask = 64'h111F111F111F111F;
defparam \Selector22~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector21~0 (
	.dataa(!logical_ch_addr[6]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~0 .extended_lut = "off";
defparam \Selector21~0 .lut_mask = 64'h111F111F111F111F;
defparam \Selector21~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!logical_ch_addr[7]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h111F111F111F111F;
defparam \Selector20~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!logical_ch_addr[8]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h111F111F111F111F;
defparam \Selector19~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!logical_ch_addr[9]),
	.datab(!\Selector2~1_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!outdata_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h111F111F111F111F;
defparam \Selector18~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!\Selector8~0_combout ),
	.datab(!outdata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'h1111111111111111;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~1 (
	.dataa(!ctrl_lock),
	.datab(!\Selector4~0_combout ),
	.datac(!\Selector12~1_combout ),
	.datad(!\WideOr5~0_combout ),
	.datae(!\WideOr17~0_combout ),
	.dataf(!\Selector16~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~1 .extended_lut = "off";
defparam \Selector16~1 .lut_mask = 64'hFFFFFFFFFFFF3BFF;
defparam \Selector16~1 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_uif (
	user_reconfig_readdata_6,
	user_reconfig_readdata_7,
	user_reconfig_readdata_10,
	user_reconfig_readdata_11,
	user_reconfig_readdata_12,
	user_reconfig_readdata_13,
	user_reconfig_readdata_14,
	user_reconfig_readdata_15,
	user_reconfig_readdata_16,
	user_reconfig_readdata_17,
	user_reconfig_readdata_18,
	user_reconfig_readdata_19,
	user_reconfig_readdata_0,
	user_reconfig_readdata_1,
	user_reconfig_readdata_2,
	user_reconfig_readdata_3,
	user_reconfig_readdata_4,
	user_reconfig_readdata_5,
	Equal1,
	user_reconfig_readdata_8,
	user_reconfig_readdata_9,
	user_reconfig_readdata_20,
	user_reconfig_readdata_21,
	user_reconfig_readdata_22,
	user_reconfig_readdata_23,
	user_reconfig_readdata_24,
	user_reconfig_readdata_25,
	user_reconfig_readdata_26,
	user_reconfig_readdata_27,
	user_reconfig_readdata_28,
	user_reconfig_readdata_29,
	user_reconfig_readdata_30,
	user_reconfig_readdata_31,
	comb,
	user_reconfig_waitrequest,
	stateSTATE_IDLE,
	ifsel_notdone_resync,
	uif_addr_offset_5,
	uif_addr_offset_4,
	uif_addr_offset_0,
	uif_addr_offset_1,
	uif_addr_offset_3,
	uif_addr_offset_2,
	Decoder3,
	Decoder31,
	Decoder32,
	rtl,
	rtl1,
	rtl2,
	rtl3,
	rtl4,
	rtl5,
	rtl6,
	rtl7,
	Decoder33,
	uif_mode_1,
	uif_mode_0,
	Decoder34,
	WideOr4,
	analog_length,
	analog_length1,
	lpbk_done,
	uif_writedata_0,
	lpbk_precdr_reg,
	lpbk_postcdr_reg,
	uif_logical_ch_addr_0,
	ph_readdata_0,
	uif_writedata_1,
	uif_logical_ch_addr_1,
	ph_readdata_1,
	uif_writedata_2,
	rtl8,
	rtl9,
	rtl10,
	uif_logical_ch_addr_2,
	ph_readdata_2,
	user_reconfig_readdata_101,
	uif_writedata_3,
	rtl11,
	rtl12,
	rtl13,
	uif_logical_ch_addr_3,
	ph_readdata_3,
	uif_writedata_4,
	rtl14,
	rtl15,
	LessThan4,
	uif_logical_ch_addr_4,
	ph_readdata_4,
	uif_writedata_5,
	rtl16,
	rtl17,
	uif_logical_ch_addr_5,
	ph_readdata_5,
	uif_writedata_6,
	rtl18,
	rtl19,
	ph_readdata_6,
	uif_logical_ch_addr_6,
	user_reconfig_readdata_71,
	rtl20,
	rtl21,
	ph_readdata_7,
	uif_logical_ch_addr_7,
	rtl22,
	Equal6,
	uif_logical_ch_addr_8,
	ph_readdata_8,
	rtl23,
	ph_readdata_9,
	uif_logical_ch_addr_9,
	uif_illegal_pch_error,
	uif_illegal_offset_error,
	ph_readdata_10,
	rtl24,
	ph_readdata_11,
	rtl25,
	ph_readdata_12,
	rtl26,
	ph_readdata_13,
	rtl27,
	ph_readdata_14,
	rtl28,
	ph_readdata_15,
	rtl29,
	ph_readdata_16,
	rtl30,
	ph_readdata_17,
	rtl31,
	ph_readdata_18,
	rtl32,
	ph_readdata_19,
	ShiftRight0,
	ph_readdata_20,
	ph_readdata_21,
	ph_readdata_22,
	ph_readdata_23,
	ph_readdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	uif_go1,
	uif_mode_01,
	Mux0,
	Mux3,
	WideOr0,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_6;
output 	user_reconfig_readdata_7;
output 	user_reconfig_readdata_10;
output 	user_reconfig_readdata_11;
output 	user_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
output 	user_reconfig_readdata_0;
output 	user_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
input 	Equal1;
output 	user_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
output 	user_reconfig_readdata_20;
output 	user_reconfig_readdata_21;
output 	user_reconfig_readdata_22;
output 	user_reconfig_readdata_23;
output 	user_reconfig_readdata_24;
output 	user_reconfig_readdata_25;
output 	user_reconfig_readdata_26;
output 	user_reconfig_readdata_27;
output 	user_reconfig_readdata_28;
output 	user_reconfig_readdata_29;
output 	user_reconfig_readdata_30;
output 	user_reconfig_readdata_31;
input 	comb;
output 	user_reconfig_waitrequest;
input 	stateSTATE_IDLE;
input 	ifsel_notdone_resync;
output 	uif_addr_offset_5;
output 	uif_addr_offset_4;
output 	uif_addr_offset_0;
output 	uif_addr_offset_1;
output 	uif_addr_offset_3;
output 	uif_addr_offset_2;
input 	Decoder3;
input 	Decoder31;
input 	Decoder32;
input 	rtl;
input 	rtl1;
input 	rtl2;
input 	rtl3;
input 	rtl4;
input 	rtl5;
input 	rtl6;
input 	rtl7;
input 	Decoder33;
output 	uif_mode_1;
output 	uif_mode_0;
input 	Decoder34;
input 	WideOr4;
input 	analog_length;
input 	analog_length1;
input 	lpbk_done;
output 	uif_writedata_0;
input 	lpbk_precdr_reg;
input 	lpbk_postcdr_reg;
output 	uif_logical_ch_addr_0;
input 	ph_readdata_0;
output 	uif_writedata_1;
output 	uif_logical_ch_addr_1;
input 	ph_readdata_1;
output 	uif_writedata_2;
input 	rtl8;
input 	rtl9;
input 	rtl10;
output 	uif_logical_ch_addr_2;
input 	ph_readdata_2;
input 	user_reconfig_readdata_101;
output 	uif_writedata_3;
input 	rtl11;
input 	rtl12;
input 	rtl13;
output 	uif_logical_ch_addr_3;
input 	ph_readdata_3;
output 	uif_writedata_4;
input 	rtl14;
input 	rtl15;
input 	LessThan4;
output 	uif_logical_ch_addr_4;
input 	ph_readdata_4;
output 	uif_writedata_5;
input 	rtl16;
input 	rtl17;
output 	uif_logical_ch_addr_5;
input 	ph_readdata_5;
output 	uif_writedata_6;
input 	rtl18;
input 	rtl19;
input 	ph_readdata_6;
output 	uif_logical_ch_addr_6;
output 	user_reconfig_readdata_71;
input 	rtl20;
input 	rtl21;
input 	ph_readdata_7;
output 	uif_logical_ch_addr_7;
input 	rtl22;
input 	Equal6;
output 	uif_logical_ch_addr_8;
input 	ph_readdata_8;
input 	rtl23;
input 	ph_readdata_9;
output 	uif_logical_ch_addr_9;
input 	uif_illegal_pch_error;
input 	uif_illegal_offset_error;
input 	ph_readdata_10;
input 	rtl24;
input 	ph_readdata_11;
input 	rtl25;
input 	ph_readdata_12;
input 	rtl26;
input 	ph_readdata_13;
input 	rtl27;
input 	ph_readdata_14;
input 	rtl28;
input 	ph_readdata_15;
input 	rtl29;
input 	ph_readdata_16;
input 	rtl30;
input 	ph_readdata_17;
input 	rtl31;
input 	ph_readdata_18;
input 	rtl32;
input 	ph_readdata_19;
input 	ShiftRight0;
input 	ph_readdata_20;
input 	ph_readdata_21;
input 	ph_readdata_22;
input 	ph_readdata_23;
input 	ph_readdata_24;
input 	ph_readdata_25;
input 	ph_readdata_26;
input 	ph_readdata_27;
input 	ph_readdata_28;
input 	ph_readdata_29;
input 	ph_readdata_30;
input 	ph_readdata_31;
output 	uif_go1;
output 	uif_mode_01;
input 	Mux0;
input 	Mux3;
output 	WideOr0;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \user_reconfig_readdata[6]~13_combout ;
wire \user_reconfig_readdata[6]~14_combout ;
wire \user_reconfig_readdata[6]~15_combout ;
wire \user_reconfig_readdata[0]~5_combout ;
wire \always0~0_combout ;
wire \uif_writedata[0]~0_combout ;
wire \uif_writedata[7]~q ;
wire \user_reconfig_readdata[7]~17_combout ;
wire \user_reconfig_readdata[7]~37_combout ;
wire \uif_writedata[10]~q ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \user_reconfig_readdata[17]~22_combout ;
wire \user_reconfig_readdata[10]~23_combout ;
wire \uif_writedata[11]~q ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \uif_writedata[12]~q ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \uif_writedata[13]~q ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \uif_writedata[14]~q ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \uif_writedata[15]~q ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \uif_writedata[16]~q ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \uif_writedata[17]~q ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \uif_writedata[18]~q ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \uif_writedata[19]~q ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \user_reconfig_readdata[0]~0_combout ;
wire \user_reconfig_readdata[0]~1_combout ;
wire \user_reconfig_readdata[0]~3_combout ;
wire \user_reconfig_readdata[0]~2_combout ;
wire \user_reconfig_readdata[0]~70_combout ;
wire \user_reconfig_readdata[0]~4_combout ;
wire \user_reconfig_readdata[0]~66_combout ;
wire \user_reconfig_readdata[1]~6_combout ;
wire \user_reconfig_readdata[1]~65_combout ;
wire \user_reconfig_readdata[1]~7_combout ;
wire \user_reconfig_readdata[1]~8_combout ;
wire \user_reconfig_readdata[1]~61_combout ;
wire \user_reconfig_readdata[2]~9_combout ;
wire \user_reconfig_readdata[2]~10_combout ;
wire \user_reconfig_readdata[2]~57_combout ;
wire \user_reconfig_readdata[3]~11_combout ;
wire \user_reconfig_readdata[3]~53_combout ;
wire \user_reconfig_readdata[4]~12_combout ;
wire \user_reconfig_readdata[4]~49_combout ;
wire \user_reconfig_readdata[5]~45_combout ;
wire \user_reconfig_readdata[5]~41_combout ;
wire \Mux27~0_combout ;
wire \user_reconfig_readdata[8]~18_combout ;
wire \user_reconfig_readdata[8]~19_combout ;
wire \uif_writedata[8]~q ;
wire \Mux27~1_combout ;
wire \Mux27~2_combout ;
wire \user_reconfig_readdata[8]~20_combout ;
wire \user_reconfig_readdata[8]~21_combout ;
wire \Mux26~0_combout ;
wire \illegal_addr_error~0_combout ;
wire \illegal_addr_error~q ;
wire \Mux26~2_combout ;
wire \uif_writedata[9]~q ;
wire \Mux26~1_combout ;
wire \user_reconfig_readdata[22]~24_combout ;
wire \user_reconfig_readdata[22]~25_combout ;
wire \Mux15~0_combout ;
wire \user_reconfig_readdata[22]~26_combout ;
wire \user_reconfig_readdata[22]~27_combout ;
wire \uif_writedata[20]~q ;
wire \Mux15~1_combout ;
wire \Mux14~0_combout ;
wire \uif_writedata[21]~q ;
wire \Mux14~1_combout ;
wire \Mux13~0_combout ;
wire \uif_writedata[22]~q ;
wire \Mux13~1_combout ;
wire \Mux12~0_combout ;
wire \uif_writedata[23]~q ;
wire \Mux12~1_combout ;
wire \user_reconfig_readdata[26]~28_combout ;
wire \user_reconfig_readdata[26]~29_combout ;
wire \user_reconfig_readdata[26]~30_combout ;
wire \user_reconfig_readdata[26]~31_combout ;
wire \user_reconfig_readdata[26]~32_combout ;
wire \uif_writedata[24]~q ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux11~2_combout ;
wire \uif_writedata[25]~q ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \uif_writedata[26]~q ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \uif_writedata[27]~q ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \user_reconfig_readdata[29]~33_combout ;
wire \user_reconfig_readdata[29]~34_combout ;
wire \user_reconfig_readdata[29]~35_combout ;
wire \user_reconfig_readdata[29]~36_combout ;
wire \uif_writedata[28]~q ;
wire \Mux7~0_combout ;
wire \uif_writedata[29]~q ;
wire \Mux6~0_combout ;
wire \uif_writedata[30]~q ;
wire \Mux5~0_combout ;
wire \uif_writedata[31]~q ;
wire \Mux4~0_combout ;
wire \uif_addr_offset[0]~0_combout ;
wire \uif_mode[1]~2_combout ;
wire \Mux0~0_combout ;
wire \uif_mode[0]~1_combout ;
wire \uif_logical_ch_addr[0]~0_combout ;
wire \Mux0~1_combout ;


RECONFIGURE_IP_altera_wait_generate wait_gen(
	.launch_signal(comb),
	.wait_req(user_reconfig_waitrequest),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.mgmt_clk_clk(mgmt_clk_clk));

dffeas \user_reconfig_readdata[6] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[6]~15_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(reconfig_mgmt_address_1),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_6),
	.prn(vcc));
defparam \user_reconfig_readdata[6] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[6] .power_up = "low";

dffeas \user_reconfig_readdata[7] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[7]~37_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(reconfig_mgmt_address_1),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_7),
	.prn(vcc));
defparam \user_reconfig_readdata[7] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[7] .power_up = "low";

dffeas \user_reconfig_readdata[10] (
	.clk(mgmt_clk_clk),
	.d(\Mux25~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_10),
	.prn(vcc));
defparam \user_reconfig_readdata[10] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[10] .power_up = "low";

dffeas \user_reconfig_readdata[11] (
	.clk(mgmt_clk_clk),
	.d(\Mux24~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_11),
	.prn(vcc));
defparam \user_reconfig_readdata[11] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[11] .power_up = "low";

dffeas \user_reconfig_readdata[12] (
	.clk(mgmt_clk_clk),
	.d(\Mux23~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_12),
	.prn(vcc));
defparam \user_reconfig_readdata[12] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[12] .power_up = "low";

dffeas \user_reconfig_readdata[13] (
	.clk(mgmt_clk_clk),
	.d(\Mux22~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_13),
	.prn(vcc));
defparam \user_reconfig_readdata[13] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[13] .power_up = "low";

dffeas \user_reconfig_readdata[14] (
	.clk(mgmt_clk_clk),
	.d(\Mux21~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_14),
	.prn(vcc));
defparam \user_reconfig_readdata[14] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[14] .power_up = "low";

dffeas \user_reconfig_readdata[15] (
	.clk(mgmt_clk_clk),
	.d(\Mux20~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_15),
	.prn(vcc));
defparam \user_reconfig_readdata[15] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[15] .power_up = "low";

dffeas \user_reconfig_readdata[16] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_16),
	.prn(vcc));
defparam \user_reconfig_readdata[16] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[16] .power_up = "low";

dffeas \user_reconfig_readdata[17] (
	.clk(mgmt_clk_clk),
	.d(\Mux18~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_17),
	.prn(vcc));
defparam \user_reconfig_readdata[17] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[17] .power_up = "low";

dffeas \user_reconfig_readdata[18] (
	.clk(mgmt_clk_clk),
	.d(\Mux17~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_18),
	.prn(vcc));
defparam \user_reconfig_readdata[18] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[18] .power_up = "low";

dffeas \user_reconfig_readdata[19] (
	.clk(mgmt_clk_clk),
	.d(\Mux16~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(\user_reconfig_readdata[17]~22_combout ),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_19),
	.prn(vcc));
defparam \user_reconfig_readdata[19] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[19] .power_up = "low";

dffeas \user_reconfig_readdata[0] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[0]~66_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_0),
	.prn(vcc));
defparam \user_reconfig_readdata[0] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[0] .power_up = "low";

dffeas \user_reconfig_readdata[1] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[1]~61_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_1),
	.prn(vcc));
defparam \user_reconfig_readdata[1] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[1] .power_up = "low";

dffeas \user_reconfig_readdata[2] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[2]~57_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_2),
	.prn(vcc));
defparam \user_reconfig_readdata[2] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[2] .power_up = "low";

dffeas \user_reconfig_readdata[3] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[3]~53_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_3),
	.prn(vcc));
defparam \user_reconfig_readdata[3] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[3] .power_up = "low";

dffeas \user_reconfig_readdata[4] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[4]~49_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_4),
	.prn(vcc));
defparam \user_reconfig_readdata[4] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[4] .power_up = "low";

dffeas \user_reconfig_readdata[5] (
	.clk(mgmt_clk_clk),
	.d(\user_reconfig_readdata[5]~41_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~5_combout ),
	.q(user_reconfig_readdata_5),
	.prn(vcc));
defparam \user_reconfig_readdata[5] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[5] .power_up = "low";

dffeas \user_reconfig_readdata[8] (
	.clk(mgmt_clk_clk),
	.d(\Mux27~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[8]~21_combout ),
	.q(user_reconfig_readdata_8),
	.prn(vcc));
defparam \user_reconfig_readdata[8] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[8] .power_up = "low";

dffeas \user_reconfig_readdata[9] (
	.clk(mgmt_clk_clk),
	.d(\Mux26~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[8]~21_combout ),
	.q(user_reconfig_readdata_9),
	.prn(vcc));
defparam \user_reconfig_readdata[9] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[9] .power_up = "low";

dffeas \user_reconfig_readdata[20] (
	.clk(mgmt_clk_clk),
	.d(\Mux15~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_20),
	.prn(vcc));
defparam \user_reconfig_readdata[20] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[20] .power_up = "low";

dffeas \user_reconfig_readdata[21] (
	.clk(mgmt_clk_clk),
	.d(\Mux14~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_21),
	.prn(vcc));
defparam \user_reconfig_readdata[21] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[21] .power_up = "low";

dffeas \user_reconfig_readdata[22] (
	.clk(mgmt_clk_clk),
	.d(\Mux13~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_22),
	.prn(vcc));
defparam \user_reconfig_readdata[22] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[22] .power_up = "low";

dffeas \user_reconfig_readdata[23] (
	.clk(mgmt_clk_clk),
	.d(\Mux12~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_23),
	.prn(vcc));
defparam \user_reconfig_readdata[23] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[23] .power_up = "low";

dffeas \user_reconfig_readdata[24] (
	.clk(mgmt_clk_clk),
	.d(\Mux11~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_24),
	.prn(vcc));
defparam \user_reconfig_readdata[24] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[24] .power_up = "low";

dffeas \user_reconfig_readdata[25] (
	.clk(mgmt_clk_clk),
	.d(\Mux10~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_25),
	.prn(vcc));
defparam \user_reconfig_readdata[25] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[25] .power_up = "low";

dffeas \user_reconfig_readdata[26] (
	.clk(mgmt_clk_clk),
	.d(\Mux9~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_26),
	.prn(vcc));
defparam \user_reconfig_readdata[26] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[26] .power_up = "low";

dffeas \user_reconfig_readdata[27] (
	.clk(mgmt_clk_clk),
	.d(\Mux8~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_27),
	.prn(vcc));
defparam \user_reconfig_readdata[27] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[27] .power_up = "low";

dffeas \user_reconfig_readdata[28] (
	.clk(mgmt_clk_clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_28),
	.prn(vcc));
defparam \user_reconfig_readdata[28] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[28] .power_up = "low";

dffeas \user_reconfig_readdata[29] (
	.clk(mgmt_clk_clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_29),
	.prn(vcc));
defparam \user_reconfig_readdata[29] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[29] .power_up = "low";

dffeas \user_reconfig_readdata[30] (
	.clk(mgmt_clk_clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_30),
	.prn(vcc));
defparam \user_reconfig_readdata[30] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[30] .power_up = "low";

dffeas \user_reconfig_readdata[31] (
	.clk(mgmt_clk_clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~23_combout ),
	.q(user_reconfig_readdata_31),
	.prn(vcc));
defparam \user_reconfig_readdata[31] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[31] .power_up = "low";

dffeas \uif_addr_offset[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_5),
	.prn(vcc));
defparam \uif_addr_offset[5] .is_wysiwyg = "true";
defparam \uif_addr_offset[5] .power_up = "low";

dffeas \uif_addr_offset[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_4),
	.prn(vcc));
defparam \uif_addr_offset[4] .is_wysiwyg = "true";
defparam \uif_addr_offset[4] .power_up = "low";

dffeas \uif_addr_offset[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_0),
	.prn(vcc));
defparam \uif_addr_offset[0] .is_wysiwyg = "true";
defparam \uif_addr_offset[0] .power_up = "low";

dffeas \uif_addr_offset[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_1),
	.prn(vcc));
defparam \uif_addr_offset[1] .is_wysiwyg = "true";
defparam \uif_addr_offset[1] .power_up = "low";

dffeas \uif_addr_offset[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_3),
	.prn(vcc));
defparam \uif_addr_offset[3] .is_wysiwyg = "true";
defparam \uif_addr_offset[3] .power_up = "low";

dffeas \uif_addr_offset[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_2),
	.prn(vcc));
defparam \uif_addr_offset[2] .is_wysiwyg = "true";
defparam \uif_addr_offset[2] .power_up = "low";

dffeas \uif_mode[1] (
	.clk(mgmt_clk_clk),
	.d(\uif_mode[1]~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_mode[0]~1_combout ),
	.q(uif_mode_1),
	.prn(vcc));
defparam \uif_mode[1] .is_wysiwyg = "true";
defparam \uif_mode[1] .power_up = "low";

dffeas \uif_mode[0] (
	.clk(mgmt_clk_clk),
	.d(Mux3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_mode[0]~1_combout ),
	.q(uif_mode_0),
	.prn(vcc));
defparam \uif_mode[0] .is_wysiwyg = "true";
defparam \uif_mode[0] .power_up = "low";

dffeas \uif_writedata[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_0),
	.prn(vcc));
defparam \uif_writedata[0] .is_wysiwyg = "true";
defparam \uif_writedata[0] .power_up = "low";

dffeas \uif_logical_ch_addr[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_0),
	.prn(vcc));
defparam \uif_logical_ch_addr[0] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[0] .power_up = "low";

dffeas \uif_writedata[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_1),
	.prn(vcc));
defparam \uif_writedata[1] .is_wysiwyg = "true";
defparam \uif_writedata[1] .power_up = "low";

dffeas \uif_logical_ch_addr[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_1),
	.prn(vcc));
defparam \uif_logical_ch_addr[1] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[1] .power_up = "low";

dffeas \uif_writedata[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_2),
	.prn(vcc));
defparam \uif_writedata[2] .is_wysiwyg = "true";
defparam \uif_writedata[2] .power_up = "low";

dffeas \uif_logical_ch_addr[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_2),
	.prn(vcc));
defparam \uif_logical_ch_addr[2] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[2] .power_up = "low";

dffeas \uif_writedata[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_3),
	.prn(vcc));
defparam \uif_writedata[3] .is_wysiwyg = "true";
defparam \uif_writedata[3] .power_up = "low";

dffeas \uif_logical_ch_addr[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_3),
	.prn(vcc));
defparam \uif_logical_ch_addr[3] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[3] .power_up = "low";

dffeas \uif_writedata[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_4),
	.prn(vcc));
defparam \uif_writedata[4] .is_wysiwyg = "true";
defparam \uif_writedata[4] .power_up = "low";

dffeas \uif_logical_ch_addr[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_4),
	.prn(vcc));
defparam \uif_logical_ch_addr[4] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[4] .power_up = "low";

dffeas \uif_writedata[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_5),
	.prn(vcc));
defparam \uif_writedata[5] .is_wysiwyg = "true";
defparam \uif_writedata[5] .power_up = "low";

dffeas \uif_logical_ch_addr[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_5),
	.prn(vcc));
defparam \uif_logical_ch_addr[5] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[5] .power_up = "low";

dffeas \uif_writedata[6] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_6),
	.prn(vcc));
defparam \uif_writedata[6] .is_wysiwyg = "true";
defparam \uif_writedata[6] .power_up = "low";

dffeas \uif_logical_ch_addr[6] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_6),
	.prn(vcc));
defparam \uif_logical_ch_addr[6] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[6] .power_up = "low";

cyclonev_lcell_comb \user_reconfig_readdata[7]~16 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(user_reconfig_readdata_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[7]~16 .extended_lut = "off";
defparam \user_reconfig_readdata[7]~16 .lut_mask = 64'h4444444444444444;
defparam \user_reconfig_readdata[7]~16 .shared_arith = "off";

dffeas \uif_logical_ch_addr[7] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_7),
	.prn(vcc));
defparam \uif_logical_ch_addr[7] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[7] .power_up = "low";

dffeas \uif_logical_ch_addr[8] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_8),
	.prn(vcc));
defparam \uif_logical_ch_addr[8] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[8] .power_up = "low";

dffeas \uif_logical_ch_addr[9] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_9),
	.prn(vcc));
defparam \uif_logical_ch_addr[9] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[9] .power_up = "low";

dffeas uif_go(
	.clk(mgmt_clk_clk),
	.d(\Mux0~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_go1),
	.prn(vcc));
defparam uif_go.is_wysiwyg = "true";
defparam uif_go.power_up = "low";

cyclonev_lcell_comb \uif_mode[0]~0 (
	.dataa(!reconfig_mgmt_writedata_0),
	.datab(!reconfig_mgmt_writedata_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(uif_mode_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_mode[0]~0 .extended_lut = "off";
defparam \uif_mode[0]~0 .lut_mask = 64'h8888888888888888;
defparam \uif_mode[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h0707070707070707;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[6]~13 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!WideOr4),
	.datad(!analog_length),
	.datae(!analog_length1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[6]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[6]~13 .extended_lut = "off";
defparam \user_reconfig_readdata[6]~13 .lut_mask = 64'h4444444C4444444C;
defparam \user_reconfig_readdata[6]~13 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[6]~14 (
	.dataa(!user_reconfig_readdata_6),
	.datab(!uif_mode_1),
	.datac(!uif_mode_0),
	.datad(!uif_writedata_6),
	.datae(!rtl19),
	.dataf(!\user_reconfig_readdata[6]~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[6]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[6]~14 .extended_lut = "off";
defparam \user_reconfig_readdata[6]~14 .lut_mask = 64'h010D010D010DF3FF;
defparam \user_reconfig_readdata[6]~14 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[6]~15 (
	.dataa(!reconfig_mgmt_address_0),
	.datab(!reconfig_mgmt_address_2),
	.datac(!\user_reconfig_readdata[6]~14_combout ),
	.datad(!ph_readdata_6),
	.datae(!uif_logical_ch_addr_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[6]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[6]~15 .extended_lut = "off";
defparam \user_reconfig_readdata[6]~15 .lut_mask = 64'h02468ACE02468ACE;
defparam \user_reconfig_readdata[6]~15 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~5 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!comb),
	.datae(!stateSTATE_IDLE),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~5 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~5 .lut_mask = 64'h00FF00D700FF00D7;
defparam \user_reconfig_readdata[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!Equal1),
	.datab(!reconfig_mgmt_write),
	.datac(!stateSTATE_IDLE),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h1010101010101010;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_writedata[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_writedata[0]~0 .extended_lut = "off";
defparam \uif_writedata[0]~0 .lut_mask = 64'h0008000800080008;
defparam \uif_writedata[0]~0 .shared_arith = "off";

dffeas \uif_writedata[7] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[7]~q ),
	.prn(vcc));
defparam \uif_writedata[7] .is_wysiwyg = "true";
defparam \uif_writedata[7] .power_up = "low";

cyclonev_lcell_comb \user_reconfig_readdata[7]~17 (
	.dataa(!user_reconfig_readdata_7),
	.datab(!uif_mode_1),
	.datac(!uif_mode_0),
	.datad(!\uif_writedata[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[7]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[7]~17 .extended_lut = "off";
defparam \user_reconfig_readdata[7]~17 .lut_mask = 64'h010D010D010D010D;
defparam \user_reconfig_readdata[7]~17 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[7]~37 (
	.dataa(!uif_logical_ch_addr_7),
	.datab(!\user_reconfig_readdata[7]~17_combout ),
	.datac(!user_reconfig_readdata_71),
	.datad(!rtl21),
	.datae(!reconfig_mgmt_address_2),
	.dataf(!reconfig_mgmt_address_0),
	.datag(!ph_readdata_7),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[7]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[7]~37 .extended_lut = "on";
defparam \user_reconfig_readdata[7]~37 .lut_mask = 64'h5555333F0F0F0000;
defparam \user_reconfig_readdata[7]~37 .shared_arith = "off";

dffeas \uif_writedata[10] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_10),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[10]~q ),
	.prn(vcc));
defparam \uif_writedata[10] .is_wysiwyg = "true";
defparam \uif_writedata[10] .power_up = "low";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!rtl8),
	.datab(!rtl18),
	.datac(!rtl9),
	.datad(!rtl24),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "off";
defparam \Mux25~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_10),
	.datad(!\uif_writedata[10]~q ),
	.datae(!\Mux25~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~1 .extended_lut = "off";
defparam \Mux25~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux25~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[17]~22 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!uif_mode_1),
	.datae(!uif_mode_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[17]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[17]~22 .extended_lut = "off";
defparam \user_reconfig_readdata[17]~22 .lut_mask = 64'hDFD7D7D7DFD7D7D7;
defparam \user_reconfig_readdata[17]~22 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[10]~23 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!comb),
	.datac(!stateSTATE_IDLE),
	.datad(!uif_mode_1),
	.datae(!uif_mode_0),
	.dataf(!user_reconfig_readdata_101),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[10]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[10]~23 .extended_lut = "off";
defparam \user_reconfig_readdata[10]~23 .lut_mask = 64'h3030302033333333;
defparam \user_reconfig_readdata[10]~23 .shared_arith = "off";

dffeas \uif_writedata[11] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_11),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[11]~q ),
	.prn(vcc));
defparam \uif_writedata[11] .is_wysiwyg = "true";
defparam \uif_writedata[11] .power_up = "low";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!rtl11),
	.datab(!rtl20),
	.datac(!rtl12),
	.datad(!rtl25),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "off";
defparam \Mux24~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_11),
	.datad(!\uif_writedata[11]~q ),
	.datae(!\Mux24~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~1 .extended_lut = "off";
defparam \Mux24~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux24~1 .shared_arith = "off";

dffeas \uif_writedata[12] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_12),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[12]~q ),
	.prn(vcc));
defparam \uif_writedata[12] .is_wysiwyg = "true";
defparam \uif_writedata[12] .power_up = "low";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!rtl1),
	.datab(!rtl22),
	.datac(!rtl14),
	.datad(!rtl26),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "off";
defparam \Mux23~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux23~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux23~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_12),
	.datad(!\uif_writedata[12]~q ),
	.datae(!\Mux23~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~1 .extended_lut = "off";
defparam \Mux23~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux23~1 .shared_arith = "off";

dffeas \uif_writedata[13] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_13),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[13]~q ),
	.prn(vcc));
defparam \uif_writedata[13] .is_wysiwyg = "true";
defparam \uif_writedata[13] .power_up = "low";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!rtl6),
	.datab(!rtl23),
	.datac(!rtl16),
	.datad(!rtl27),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "off";
defparam \Mux22~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux22~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux22~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_13),
	.datad(!\uif_writedata[13]~q ),
	.datae(!\Mux22~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~1 .extended_lut = "off";
defparam \Mux22~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux22~1 .shared_arith = "off";

dffeas \uif_writedata[14] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_14),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[14]~q ),
	.prn(vcc));
defparam \uif_writedata[14] .is_wysiwyg = "true";
defparam \uif_writedata[14] .power_up = "low";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!rtl9),
	.datab(!rtl24),
	.datac(!rtl18),
	.datad(!rtl28),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "off";
defparam \Mux21~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux21~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_14),
	.datad(!\uif_writedata[14]~q ),
	.datae(!\Mux21~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~1 .extended_lut = "off";
defparam \Mux21~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux21~1 .shared_arith = "off";

dffeas \uif_writedata[15] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_15),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[15]~q ),
	.prn(vcc));
defparam \uif_writedata[15] .is_wysiwyg = "true";
defparam \uif_writedata[15] .power_up = "low";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!rtl12),
	.datab(!rtl25),
	.datac(!rtl20),
	.datad(!rtl29),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "off";
defparam \Mux20~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux20~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_15),
	.datad(!\uif_writedata[15]~q ),
	.datae(!\Mux20~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~1 .extended_lut = "off";
defparam \Mux20~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux20~1 .shared_arith = "off";

dffeas \uif_writedata[16] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_16),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[16]~q ),
	.prn(vcc));
defparam \uif_writedata[16] .is_wysiwyg = "true";
defparam \uif_writedata[16] .power_up = "low";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!rtl14),
	.datab(!rtl26),
	.datac(!rtl22),
	.datad(!rtl30),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "off";
defparam \Mux19~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux19~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_16),
	.datad(!\uif_writedata[16]~q ),
	.datae(!\Mux19~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~1 .extended_lut = "off";
defparam \Mux19~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux19~1 .shared_arith = "off";

dffeas \uif_writedata[17] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_17),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[17]~q ),
	.prn(vcc));
defparam \uif_writedata[17] .is_wysiwyg = "true";
defparam \uif_writedata[17] .power_up = "low";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!rtl16),
	.datab(!rtl27),
	.datac(!rtl23),
	.datad(!rtl31),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "off";
defparam \Mux18~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux18~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux18~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_17),
	.datad(!\uif_writedata[17]~q ),
	.datae(!\Mux18~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux18~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~1 .extended_lut = "off";
defparam \Mux18~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux18~1 .shared_arith = "off";

dffeas \uif_writedata[18] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_18),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[18]~q ),
	.prn(vcc));
defparam \uif_writedata[18] .is_wysiwyg = "true";
defparam \uif_writedata[18] .power_up = "low";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!rtl18),
	.datab(!rtl28),
	.datac(!rtl24),
	.datad(!rtl32),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "off";
defparam \Mux17~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux17~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux17~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_18),
	.datad(!\uif_writedata[18]~q ),
	.datae(!\Mux17~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~1 .extended_lut = "off";
defparam \Mux17~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux17~1 .shared_arith = "off";

dffeas \uif_writedata[19] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_19),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[19]~q ),
	.prn(vcc));
defparam \uif_writedata[19] .is_wysiwyg = "true";
defparam \uif_writedata[19] .power_up = "low";

cyclonev_lcell_comb \Mux16~0 (
	.dataa(!rtl20),
	.datab(!rtl29),
	.datac(!rtl25),
	.datad(!ShiftRight0),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "off";
defparam \Mux16~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux16~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~1 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!ph_readdata_19),
	.datad(!\uif_writedata[19]~q ),
	.datae(!\Mux16~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~1 .extended_lut = "off";
defparam \Mux16~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux16~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~0 (
	.dataa(!Decoder33),
	.datab(!uif_mode_1),
	.datac(!uif_mode_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~0 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~0 .lut_mask = 64'h8080808080808080;
defparam \user_reconfig_readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~1 (
	.dataa(!Decoder32),
	.datab(!\user_reconfig_readdata[0]~0_combout ),
	.datac(!Decoder34),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~1 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~1 .lut_mask = 64'h0202020202020202;
defparam \user_reconfig_readdata[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~3 (
	.dataa(!lpbk_precdr_reg),
	.datab(!Decoder32),
	.datac(!\user_reconfig_readdata[0]~0_combout ),
	.datad(!lpbk_postcdr_reg),
	.datae(!Decoder3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~3 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~3 .lut_mask = 64'h0101010D0101010D;
defparam \user_reconfig_readdata[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~2 (
	.dataa(!Decoder33),
	.datab(!WideOr4),
	.datac(!analog_length),
	.datad(!analog_length1),
	.datae(!lpbk_done),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~2 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~2 .lut_mask = 64'h55557FFF55557FFF;
defparam \user_reconfig_readdata[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~70 (
	.dataa(!\user_reconfig_readdata[0]~3_combout ),
	.datab(!uif_writedata_0),
	.datac(!user_reconfig_readdata_0),
	.datad(!\user_reconfig_readdata[0]~2_combout ),
	.datae(!uif_mode_0),
	.dataf(!uif_mode_1),
	.datag(!rtl4),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~70 .extended_lut = "on";
defparam \user_reconfig_readdata[0]~70 .lut_mask = 64'h555F77775F5F5F5F;
defparam \user_reconfig_readdata[0]~70 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~4 (
	.dataa(!Decoder3),
	.datab(!rtl4),
	.datac(!rtl7),
	.datad(!\user_reconfig_readdata[0]~1_combout ),
	.datae(!\user_reconfig_readdata[0]~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~4 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~4 .lut_mask = 64'h0008FFFF0008FFFF;
defparam \user_reconfig_readdata[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~66 (
	.dataa(!ph_readdata_0),
	.datab(!uif_logical_ch_addr_0),
	.datac(!\user_reconfig_readdata[0]~4_combout ),
	.datad(!reconfig_mgmt_address_0),
	.datae(!reconfig_mgmt_address_2),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_addr_offset_0),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~66 .extended_lut = "on";
defparam \user_reconfig_readdata[0]~66 .lut_mask = 64'h33550F00000F0000;
defparam \user_reconfig_readdata[0]~66 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[1]~6 (
	.dataa(!Decoder34),
	.datab(!rtl4),
	.datac(!analog_length),
	.datad(!analog_length1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[1]~6 .extended_lut = "off";
defparam \user_reconfig_readdata[1]~6 .lut_mask = 64'hE444E444E444E444;
defparam \user_reconfig_readdata[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[1]~65 (
	.dataa(!uif_addr_offset_5),
	.datab(!uif_addr_offset_4),
	.datac(!uif_addr_offset_1),
	.datad(!uif_addr_offset_0),
	.datae(!uif_mode_0),
	.dataf(!Decoder31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[1]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[1]~65 .extended_lut = "off";
defparam \user_reconfig_readdata[1]~65 .lut_mask = 64'hFFFF00009FFF0000;
defparam \user_reconfig_readdata[1]~65 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[1]~7 (
	.dataa(!user_reconfig_readdata_1),
	.datab(!uif_mode_1),
	.datac(!uif_mode_0),
	.datad(!rtl7),
	.datae(!uif_writedata_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[1]~7 .extended_lut = "off";
defparam \user_reconfig_readdata[1]~7 .lut_mask = 64'h01310D3D01310D3D;
defparam \user_reconfig_readdata[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[1]~8 (
	.dataa(!Decoder3),
	.datab(!rtl7),
	.datac(!\user_reconfig_readdata[1]~6_combout ),
	.datad(!\user_reconfig_readdata[1]~65_combout ),
	.datae(!\user_reconfig_readdata[1]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[1]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[1]~8 .extended_lut = "off";
defparam \user_reconfig_readdata[1]~8 .lut_mask = 64'h0020FFFF0020FFFF;
defparam \user_reconfig_readdata[1]~8 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[1]~61 (
	.dataa(!ph_readdata_1),
	.datab(!uif_logical_ch_addr_1),
	.datac(!\user_reconfig_readdata[1]~8_combout ),
	.datad(!reconfig_mgmt_address_0),
	.datae(!reconfig_mgmt_address_2),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_addr_offset_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[1]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[1]~61 .extended_lut = "on";
defparam \user_reconfig_readdata[1]~61 .lut_mask = 64'h33550F00000F0000;
defparam \user_reconfig_readdata[1]~61 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[2]~9 (
	.dataa(!Decoder33),
	.datab(!WideOr4),
	.datac(!analog_length),
	.datad(!analog_length1),
	.datae(!lpbk_done),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[2]~9 .extended_lut = "off";
defparam \user_reconfig_readdata[2]~9 .lut_mask = 64'h00000A2A00000A2A;
defparam \user_reconfig_readdata[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[2]~10 (
	.dataa(!user_reconfig_readdata_2),
	.datab(!uif_mode_1),
	.datac(!uif_mode_0),
	.datad(!uif_writedata_2),
	.datae(!rtl10),
	.dataf(!\user_reconfig_readdata[2]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[2]~10 .extended_lut = "off";
defparam \user_reconfig_readdata[2]~10 .lut_mask = 64'h010D313D010DF1FD;
defparam \user_reconfig_readdata[2]~10 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[2]~57 (
	.dataa(!ph_readdata_2),
	.datab(!uif_logical_ch_addr_2),
	.datac(!\user_reconfig_readdata[2]~10_combout ),
	.datad(!reconfig_mgmt_address_0),
	.datae(!reconfig_mgmt_address_2),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_addr_offset_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[2]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[2]~57 .extended_lut = "on";
defparam \user_reconfig_readdata[2]~57 .lut_mask = 64'h33550F00000F0000;
defparam \user_reconfig_readdata[2]~57 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[3]~11 (
	.dataa(!user_reconfig_readdata_3),
	.datab(!uif_mode_1),
	.datac(!uif_mode_0),
	.datad(!analog_length),
	.datae(!uif_writedata_3),
	.dataf(!rtl13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[3]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[3]~11 .extended_lut = "off";
defparam \user_reconfig_readdata[3]~11 .lut_mask = 64'h01010D0D31F13DFD;
defparam \user_reconfig_readdata[3]~11 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[3]~53 (
	.dataa(!ph_readdata_3),
	.datab(!uif_logical_ch_addr_3),
	.datac(!\user_reconfig_readdata[3]~11_combout ),
	.datad(!reconfig_mgmt_address_0),
	.datae(!reconfig_mgmt_address_2),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_addr_offset_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[3]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[3]~53 .extended_lut = "on";
defparam \user_reconfig_readdata[3]~53 .lut_mask = 64'h33550F00000F0000;
defparam \user_reconfig_readdata[3]~53 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[4]~12 (
	.dataa(!user_reconfig_readdata_4),
	.datab(!uif_mode_1),
	.datac(!uif_mode_0),
	.datad(!uif_writedata_4),
	.datae(!rtl15),
	.dataf(!LessThan4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[4]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[4]~12 .extended_lut = "off";
defparam \user_reconfig_readdata[4]~12 .lut_mask = 64'h010D313D010DF1FD;
defparam \user_reconfig_readdata[4]~12 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[4]~49 (
	.dataa(!ph_readdata_4),
	.datab(!uif_logical_ch_addr_4),
	.datac(!\user_reconfig_readdata[4]~12_combout ),
	.datad(!reconfig_mgmt_address_0),
	.datae(!reconfig_mgmt_address_2),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_addr_offset_4),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[4]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[4]~49 .extended_lut = "on";
defparam \user_reconfig_readdata[4]~49 .lut_mask = 64'h33550F00000F0000;
defparam \user_reconfig_readdata[4]~49 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[5]~45 (
	.dataa(!rtl17),
	.datab(!analog_length1),
	.datac(!uif_writedata_5),
	.datad(!uif_mode_1),
	.datae(!uif_mode_0),
	.dataf(!user_reconfig_readdata_5),
	.datag(!analog_length),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[5]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[5]~45 .extended_lut = "on";
defparam \user_reconfig_readdata[5]~45 .lut_mask = 64'h01550F0001550FFF;
defparam \user_reconfig_readdata[5]~45 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[5]~41 (
	.dataa(!ph_readdata_5),
	.datab(!uif_logical_ch_addr_5),
	.datac(!\user_reconfig_readdata[5]~45_combout ),
	.datad(!reconfig_mgmt_address_0),
	.datae(!reconfig_mgmt_address_2),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_addr_offset_5),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[5]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[5]~41 .extended_lut = "on";
defparam \user_reconfig_readdata[5]~41 .lut_mask = 64'h33550F00000F0000;
defparam \user_reconfig_readdata[5]~41 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!rtl),
	.datab(!rtl14),
	.datac(!rtl1),
	.datad(!rtl22),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "off";
defparam \Mux27~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[8]~18 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!uif_mode_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[8]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[8]~18 .extended_lut = "off";
defparam \user_reconfig_readdata[8]~18 .lut_mask = 64'h0F070F070F070F07;
defparam \user_reconfig_readdata[8]~18 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[8]~19 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[8]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[8]~19 .extended_lut = "off";
defparam \user_reconfig_readdata[8]~19 .lut_mask = 64'h0F070F070F070F07;
defparam \user_reconfig_readdata[8]~19 .shared_arith = "off";

dffeas \uif_writedata[8] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[8]~q ),
	.prn(vcc));
defparam \uif_writedata[8] .is_wysiwyg = "true";
defparam \uif_writedata[8] .power_up = "low";

cyclonev_lcell_comb \Mux27~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!stateSTATE_IDLE),
	.datad(!uif_logical_ch_addr_8),
	.datae(!ph_readdata_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~1 .extended_lut = "off";
defparam \Mux27~1 .lut_mask = 64'h048C26AE048C26AE;
defparam \Mux27~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~2 (
	.dataa(!\Mux27~0_combout ),
	.datab(!\user_reconfig_readdata[8]~18_combout ),
	.datac(!\user_reconfig_readdata[8]~19_combout ),
	.datad(!\uif_writedata[8]~q ),
	.datae(!\Mux27~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~2 .extended_lut = "off";
defparam \Mux27~2 .lut_mask = 64'h0434C4F40434C4F4;
defparam \Mux27~2 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[8]~20 (
	.dataa(!reconfig_mgmt_address_0),
	.datab(!stateSTATE_IDLE),
	.datac(!uif_mode_1),
	.datad(!uif_mode_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[8]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[8]~20 .extended_lut = "off";
defparam \user_reconfig_readdata[8]~20 .lut_mask = 64'hCCC4CCC4CCC4CCC4;
defparam \user_reconfig_readdata[8]~20 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[8]~21 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!comb),
	.datae(!\user_reconfig_readdata[8]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[8]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[8]~21 .extended_lut = "off";
defparam \user_reconfig_readdata[8]~21 .lut_mask = 64'h00D700FF00D700FF;
defparam \user_reconfig_readdata[8]~21 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!rtl5),
	.datab(!rtl16),
	.datac(!rtl6),
	.datad(!rtl23),
	.datae(!rtl2),
	.dataf(!rtl3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "off";
defparam \Mux26~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \illegal_addr_error~0 (
	.dataa(!Equal1),
	.datab(!reconfig_mgmt_read),
	.datac(!reconfig_mgmt_write),
	.datad(!\illegal_addr_error~q ),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\illegal_addr_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \illegal_addr_error~0 .extended_lut = "off";
defparam \illegal_addr_error~0 .lut_mask = 64'h000015FF000015FF;
defparam \illegal_addr_error~0 .shared_arith = "off";

dffeas illegal_addr_error(
	.clk(mgmt_clk_clk),
	.d(\illegal_addr_error~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\illegal_addr_error~q ),
	.prn(vcc));
defparam illegal_addr_error.is_wysiwyg = "true";
defparam illegal_addr_error.power_up = "low";

cyclonev_lcell_comb \Mux26~2 (
	.dataa(!uif_illegal_offset_error),
	.datab(!uif_illegal_pch_error),
	.datac(!ph_readdata_9),
	.datad(!\illegal_addr_error~q ),
	.datae(!reconfig_mgmt_address_0),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_logical_ch_addr_9),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~2 .extended_lut = "on";
defparam \Mux26~2 .lut_mask = 64'h0F0F0F0F77FF0000;
defparam \Mux26~2 .shared_arith = "off";

dffeas \uif_writedata[9] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[9]~q ),
	.prn(vcc));
defparam \uif_writedata[9] .is_wysiwyg = "true";
defparam \uif_writedata[9] .power_up = "low";

cyclonev_lcell_comb \Mux26~1 (
	.dataa(!\user_reconfig_readdata[8]~18_combout ),
	.datab(!\user_reconfig_readdata[8]~19_combout ),
	.datac(!\Mux26~0_combout ),
	.datad(!\Mux26~2_combout ),
	.datae(!\uif_writedata[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~1 .extended_lut = "off";
defparam \Mux26~1 .lut_mask = 64'h028A46CE028A46CE;
defparam \Mux26~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[22]~24 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!rtl2),
	.datad(!rtl3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[22]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[22]~24 .extended_lut = "off";
defparam \user_reconfig_readdata[22]~24 .lut_mask = 64'h0772077207720772;
defparam \user_reconfig_readdata[22]~24 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[22]~25 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!rtl2),
	.datad(!rtl3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[22]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[22]~25 .extended_lut = "off";
defparam \user_reconfig_readdata[22]~25 .lut_mask = 64'h7072707270727072;
defparam \user_reconfig_readdata[22]~25 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~0 (
	.dataa(!rtl22),
	.datab(!rtl26),
	.datac(!rtl30),
	.datad(!\user_reconfig_readdata[22]~24_combout ),
	.datae(!\user_reconfig_readdata[22]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~0 .extended_lut = "off";
defparam \Mux15~0 .lut_mask = 64'h000F5533000F5533;
defparam \Mux15~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[22]~26 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!user_reconfig_readdata_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[22]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[22]~26 .extended_lut = "off";
defparam \user_reconfig_readdata[22]~26 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \user_reconfig_readdata[22]~26 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[22]~27 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[22]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[22]~27 .extended_lut = "off";
defparam \user_reconfig_readdata[22]~27 .lut_mask = 64'h2028202820282028;
defparam \user_reconfig_readdata[22]~27 .shared_arith = "off";

dffeas \uif_writedata[20] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_20),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[20]~q ),
	.prn(vcc));
defparam \uif_writedata[20] .is_wysiwyg = "true";
defparam \uif_writedata[20] .power_up = "low";

cyclonev_lcell_comb \Mux15~1 (
	.dataa(!\Mux15~0_combout ),
	.datab(!\user_reconfig_readdata[22]~26_combout ),
	.datac(!\user_reconfig_readdata[22]~27_combout ),
	.datad(!ph_readdata_20),
	.datae(!\uif_writedata[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~1 .extended_lut = "off";
defparam \Mux15~1 .lut_mask = 64'h10131C1F10131C1F;
defparam \Mux15~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!rtl23),
	.datab(!rtl27),
	.datac(!rtl31),
	.datad(!\user_reconfig_readdata[22]~24_combout ),
	.datae(!\user_reconfig_readdata[22]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "off";
defparam \Mux14~0 .lut_mask = 64'h000F5533000F5533;
defparam \Mux14~0 .shared_arith = "off";

dffeas \uif_writedata[21] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_21),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[21]~q ),
	.prn(vcc));
defparam \uif_writedata[21] .is_wysiwyg = "true";
defparam \uif_writedata[21] .power_up = "low";

cyclonev_lcell_comb \Mux14~1 (
	.dataa(!\user_reconfig_readdata[22]~26_combout ),
	.datab(!\user_reconfig_readdata[22]~27_combout ),
	.datac(!\Mux14~0_combout ),
	.datad(!ph_readdata_21),
	.datae(!\uif_writedata[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~1 .extended_lut = "off";
defparam \Mux14~1 .lut_mask = 64'h0415263704152637;
defparam \Mux14~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~0 (
	.dataa(!rtl24),
	.datab(!rtl28),
	.datac(!rtl32),
	.datad(!\user_reconfig_readdata[22]~24_combout ),
	.datae(!\user_reconfig_readdata[22]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "off";
defparam \Mux13~0 .lut_mask = 64'h000F5533000F5533;
defparam \Mux13~0 .shared_arith = "off";

dffeas \uif_writedata[22] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_22),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[22]~q ),
	.prn(vcc));
defparam \uif_writedata[22] .is_wysiwyg = "true";
defparam \uif_writedata[22] .power_up = "low";

cyclonev_lcell_comb \Mux13~1 (
	.dataa(!\user_reconfig_readdata[22]~26_combout ),
	.datab(!\user_reconfig_readdata[22]~27_combout ),
	.datac(!\Mux13~0_combout ),
	.datad(!ph_readdata_22),
	.datae(!\uif_writedata[22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~1 .extended_lut = "off";
defparam \Mux13~1 .lut_mask = 64'h0415263704152637;
defparam \Mux13~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~0 (
	.dataa(!rtl25),
	.datab(!rtl29),
	.datac(!ShiftRight0),
	.datad(!\user_reconfig_readdata[22]~24_combout ),
	.datae(!\user_reconfig_readdata[22]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "off";
defparam \Mux12~0 .lut_mask = 64'h000F5533000F5533;
defparam \Mux12~0 .shared_arith = "off";

dffeas \uif_writedata[23] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_23),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[23]~q ),
	.prn(vcc));
defparam \uif_writedata[23] .is_wysiwyg = "true";
defparam \uif_writedata[23] .power_up = "low";

cyclonev_lcell_comb \Mux12~1 (
	.dataa(!\user_reconfig_readdata[22]~26_combout ),
	.datab(!\user_reconfig_readdata[22]~27_combout ),
	.datac(!\Mux12~0_combout ),
	.datad(!ph_readdata_23),
	.datae(!\uif_writedata[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~1 .extended_lut = "off";
defparam \Mux12~1 .lut_mask = 64'h0415263704152637;
defparam \Mux12~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[26]~28 (
	.dataa(!reconfig_mgmt_address_0),
	.datab(!reconfig_mgmt_address_2),
	.datac(!uif_mode_1),
	.datad(!uif_mode_0),
	.datae(!rtl2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[26]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[26]~28 .extended_lut = "off";
defparam \user_reconfig_readdata[26]~28 .lut_mask = 64'h4666446446664464;
defparam \user_reconfig_readdata[26]~28 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[26]~29 (
	.dataa(!Equal6),
	.datab(!rtl3),
	.datac(!\user_reconfig_readdata[26]~28_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[26]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[26]~29 .extended_lut = "off";
defparam \user_reconfig_readdata[26]~29 .lut_mask = 64'h0202020202020202;
defparam \user_reconfig_readdata[26]~29 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[26]~30 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\user_reconfig_readdata[26]~29_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[26]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[26]~30 .extended_lut = "off";
defparam \user_reconfig_readdata[26]~30 .lut_mask = 64'hAA20AA20AA20AA20;
defparam \user_reconfig_readdata[26]~30 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[26]~31 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\user_reconfig_readdata[26]~29_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[26]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[26]~31 .extended_lut = "off";
defparam \user_reconfig_readdata[26]~31 .lut_mask = 64'h20AA20AA20AA20AA;
defparam \user_reconfig_readdata[26]~31 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[26]~32 (
	.dataa(!Equal6),
	.datab(!rtl3),
	.datac(!\user_reconfig_readdata[26]~28_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[26]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[26]~32 .extended_lut = "off";
defparam \user_reconfig_readdata[26]~32 .lut_mask = 64'h0707070707070707;
defparam \user_reconfig_readdata[26]~32 .shared_arith = "off";

dffeas \uif_writedata[24] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_24),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[24]~q ),
	.prn(vcc));
defparam \uif_writedata[24] .is_wysiwyg = "true";
defparam \uif_writedata[24] .power_up = "low";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!Equal6),
	.datab(!rtl3),
	.datac(!\user_reconfig_readdata[26]~28_combout ),
	.datad(!\user_reconfig_readdata[26]~31_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "off";
defparam \Mux11~0 .lut_mask = 64'h0D000D000D000D00;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~1 (
	.dataa(!rtl26),
	.datab(!\user_reconfig_readdata[26]~32_combout ),
	.datac(!\uif_writedata[24]~q ),
	.datad(!\Mux11~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~1 .extended_lut = "off";
defparam \Mux11~1 .lut_mask = 64'h0047004700470047;
defparam \Mux11~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~2 (
	.dataa(!rtl30),
	.datab(!\user_reconfig_readdata[26]~30_combout ),
	.datac(!\user_reconfig_readdata[26]~31_combout ),
	.datad(!ph_readdata_24),
	.datae(!\Mux11~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~2 .extended_lut = "off";
defparam \Mux11~2 .lut_mask = 64'h0407373704073737;
defparam \Mux11~2 .shared_arith = "off";

dffeas \uif_writedata[25] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_25),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[25]~q ),
	.prn(vcc));
defparam \uif_writedata[25] .is_wysiwyg = "true";
defparam \uif_writedata[25] .power_up = "low";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!rtl27),
	.datab(!\user_reconfig_readdata[26]~32_combout ),
	.datac(!\Mux11~0_combout ),
	.datad(!\uif_writedata[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h0407040704070407;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~1 (
	.dataa(!rtl31),
	.datab(!\user_reconfig_readdata[26]~30_combout ),
	.datac(!\user_reconfig_readdata[26]~31_combout ),
	.datad(!ph_readdata_25),
	.datae(!\Mux10~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~1 .extended_lut = "off";
defparam \Mux10~1 .lut_mask = 64'h0407373704073737;
defparam \Mux10~1 .shared_arith = "off";

dffeas \uif_writedata[26] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_26),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[26]~q ),
	.prn(vcc));
defparam \uif_writedata[26] .is_wysiwyg = "true";
defparam \uif_writedata[26] .power_up = "low";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!rtl28),
	.datab(!\user_reconfig_readdata[26]~32_combout ),
	.datac(!\Mux11~0_combout ),
	.datad(!\uif_writedata[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h0407040704070407;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~1 (
	.dataa(!rtl32),
	.datab(!\user_reconfig_readdata[26]~30_combout ),
	.datac(!\user_reconfig_readdata[26]~31_combout ),
	.datad(!ph_readdata_26),
	.datae(!\Mux9~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~1 .extended_lut = "off";
defparam \Mux9~1 .lut_mask = 64'h0407373704073737;
defparam \Mux9~1 .shared_arith = "off";

dffeas \uif_writedata[27] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_27),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[27]~q ),
	.prn(vcc));
defparam \uif_writedata[27] .is_wysiwyg = "true";
defparam \uif_writedata[27] .power_up = "low";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!rtl29),
	.datab(!\user_reconfig_readdata[26]~32_combout ),
	.datac(!\Mux11~0_combout ),
	.datad(!\uif_writedata[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h0407040704070407;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~1 (
	.dataa(!ShiftRight0),
	.datab(!\user_reconfig_readdata[26]~30_combout ),
	.datac(!\user_reconfig_readdata[26]~31_combout ),
	.datad(!ph_readdata_27),
	.datae(!\Mux8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~1 .extended_lut = "off";
defparam \Mux8~1 .lut_mask = 64'h0407373704073737;
defparam \Mux8~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[29]~33 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!rtl2),
	.datad(!rtl3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[29]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[29]~33 .extended_lut = "off";
defparam \user_reconfig_readdata[29]~33 .lut_mask = 64'h7222722272227222;
defparam \user_reconfig_readdata[29]~33 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[29]~34 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\user_reconfig_readdata[29]~33_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[29]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[29]~34 .extended_lut = "off";
defparam \user_reconfig_readdata[29]~34 .lut_mask = 64'h2028202820282028;
defparam \user_reconfig_readdata[29]~34 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[29]~35 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!\user_reconfig_readdata[29]~34_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[29]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[29]~35 .extended_lut = "off";
defparam \user_reconfig_readdata[29]~35 .lut_mask = 64'h0B0B0B0B0B0B0B0B;
defparam \user_reconfig_readdata[29]~35 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[29]~36 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal6),
	.datac(!\user_reconfig_readdata[29]~34_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[29]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[29]~36 .extended_lut = "off";
defparam \user_reconfig_readdata[29]~36 .lut_mask = 64'h0E0E0E0E0E0E0E0E;
defparam \user_reconfig_readdata[29]~36 .shared_arith = "off";

dffeas \uif_writedata[28] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_28),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[28]~q ),
	.prn(vcc));
defparam \uif_writedata[28] .is_wysiwyg = "true";
defparam \uif_writedata[28] .power_up = "low";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!rtl30),
	.datab(!\user_reconfig_readdata[29]~35_combout ),
	.datac(!\user_reconfig_readdata[29]~36_combout ),
	.datad(!ph_readdata_28),
	.datae(!\uif_writedata[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h0407343704073437;
defparam \Mux7~0 .shared_arith = "off";

dffeas \uif_writedata[29] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_29),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[29]~q ),
	.prn(vcc));
defparam \uif_writedata[29] .is_wysiwyg = "true";
defparam \uif_writedata[29] .power_up = "low";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!rtl31),
	.datab(!\user_reconfig_readdata[29]~35_combout ),
	.datac(!\user_reconfig_readdata[29]~36_combout ),
	.datad(!ph_readdata_29),
	.datae(!\uif_writedata[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h0407343704073437;
defparam \Mux6~0 .shared_arith = "off";

dffeas \uif_writedata[30] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_30),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[30]~q ),
	.prn(vcc));
defparam \uif_writedata[30] .is_wysiwyg = "true";
defparam \uif_writedata[30] .power_up = "low";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!rtl32),
	.datab(!\user_reconfig_readdata[29]~35_combout ),
	.datac(!\user_reconfig_readdata[29]~36_combout ),
	.datad(!ph_readdata_30),
	.datae(!\uif_writedata[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'h0407343704073437;
defparam \Mux5~0 .shared_arith = "off";

dffeas \uif_writedata[31] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_31),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[31]~q ),
	.prn(vcc));
defparam \uif_writedata[31] .is_wysiwyg = "true";
defparam \uif_writedata[31] .power_up = "low";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!ShiftRight0),
	.datab(!\user_reconfig_readdata[29]~35_combout ),
	.datac(!\user_reconfig_readdata[29]~36_combout ),
	.datad(!ph_readdata_31),
	.datae(!\uif_writedata[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'h0407343704073437;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_addr_offset[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_addr_offset[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_addr_offset[0]~0 .extended_lut = "off";
defparam \uif_addr_offset[0]~0 .lut_mask = 64'h0010001000100010;
defparam \uif_addr_offset[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_mode[1]~2 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_mode[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_mode[1]~2 .extended_lut = "off";
defparam \uif_mode[1]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \uif_mode[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!comb),
	.datab(!stateSTATE_IDLE),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h4444444444444444;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_mode[0]~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!\always0~0_combout ),
	.datac(!uif_mode_01),
	.datad(!\Mux0~0_combout ),
	.datae(!Mux0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_mode[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_mode[0]~1 .extended_lut = "off";
defparam \uif_mode[0]~1 .lut_mask = 64'h000010BA000010BA;
defparam \uif_mode[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \uif_logical_ch_addr[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_logical_ch_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_logical_ch_addr[0]~0 .extended_lut = "off";
defparam \uif_logical_ch_addr[0]~0 .lut_mask = 64'h0080008000800080;
defparam \uif_logical_ch_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!\always0~0_combout ),
	.datac(!uif_mode_01),
	.datad(!\Mux0~0_combout ),
	.datae(!Mux0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~1 .extended_lut = "off";
defparam \Mux0~1 .lut_mask = 64'h000010BA000010BA;
defparam \Mux0~1 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_altera_wait_generate (
	launch_signal,
	wait_req,
	ifsel_notdone_resync,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	launch_signal;
output 	wait_req;
input 	ifsel_notdone_resync;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rst_sync|resync_chains[0].sync_r[1]~q ;
wire \launch_reg~q ;
wire \wait_reg~0_combout ;
wire \wait_reg~q ;


RECONFIGURE_IP_alt_xcvr_resync rst_sync(
	.resync_chains0sync_r_1(\rst_sync|resync_chains[0].sync_r[1]~q ),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.clk(mgmt_clk_clk));

cyclonev_lcell_comb \wait_req~0 (
	.dataa(!\rst_sync|resync_chains[0].sync_r[1]~q ),
	.datab(!launch_signal),
	.datac(!\launch_reg~q ),
	.datad(!\wait_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wait_req),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_req~0 .extended_lut = "off";
defparam \wait_req~0 .lut_mask = 64'h4544454445444544;
defparam \wait_req~0 .shared_arith = "off";

dffeas launch_reg(
	.clk(mgmt_clk_clk),
	.d(launch_signal),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\launch_reg~q ),
	.prn(vcc));
defparam launch_reg.is_wysiwyg = "true";
defparam launch_reg.power_up = "low";

cyclonev_lcell_comb \wait_reg~0 (
	.dataa(!launch_signal),
	.datab(!wait_req),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_reg~0 .extended_lut = "off";
defparam \wait_reg~0 .lut_mask = 64'h1111111111111111;
defparam \wait_reg~0 .shared_arith = "off";

dffeas wait_reg(
	.clk(mgmt_clk_clk),
	.d(\wait_reg~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_reg~q ),
	.prn(vcc));
defparam wait_reg.is_wysiwyg = "true";
defparam wait_reg.power_up = "low";

endmodule

module RECONFIGURE_IP_alt_xcvr_resync (
	resync_chains0sync_r_1,
	ifsel_notdone_resync,
	clk)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
input 	ifsel_notdone_resync;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \resync_chains[0].sync_r[0]~q ;


dffeas \resync_chains[0].sync_r[1] (
	.clk(clk),
	.d(\resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resync_chains0sync_r_1),
	.prn(vcc));
defparam \resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[1] .power_up = "low";

dffeas \resync_chains[0].sync_r[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[0] .power_up = "low";

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_basic (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	Equal2,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	mutex_grant,
	master_write,
	wbasic_write_8,
	wbasic_write_81,
	wbasic_write_82,
	mutex_grant1,
	wbasic_address_2_8,
	mutex_grant2,
	wbasic_address_0_8,
	wbasic_address_1_8,
	lif_waitrequest,
	wbasic_read_8,
	wbasic_read_81,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	resync_chains0sync_r_1,
	native_reconfig_writedata_0,
	native_reconfig_writedata_1,
	native_reconfig_writedata_2,
	native_reconfig_writedata_3,
	native_reconfig_writedata_4,
	native_reconfig_writedata_5,
	native_reconfig_writedata_6,
	native_reconfig_writedata_7,
	native_reconfig_writedata_8,
	native_reconfig_writedata_9,
	native_reconfig_writedata_10,
	native_reconfig_writedata_11,
	native_reconfig_writedata_12,
	native_reconfig_writedata_13,
	native_reconfig_writedata_14,
	native_reconfig_writedata_15,
	native_reconfig_write_0,
	native_reconfig_read_0,
	native_reconfig_address_0,
	native_reconfig_address_1,
	native_reconfig_address_2,
	native_reconfig_address_3,
	native_reconfig_address_4,
	native_reconfig_address_5,
	native_reconfig_address_6,
	native_reconfig_address_7,
	native_reconfig_address_8,
	native_reconfig_address_9,
	native_reconfig_address_10,
	native_reconfig_address_11,
	pif_testbus_sel_0,
	pif_testbus_sel_1,
	pif_testbus_sel_2,
	pif_testbus_sel_3,
	pif_interface_sel,
	pif_ser_shift_load,
	native_reconfig_writedata_16,
	native_reconfig_writedata_17,
	native_reconfig_writedata_18,
	native_reconfig_writedata_19,
	native_reconfig_writedata_20,
	native_reconfig_writedata_21,
	native_reconfig_writedata_22,
	native_reconfig_writedata_23,
	native_reconfig_writedata_24,
	native_reconfig_writedata_25,
	native_reconfig_writedata_26,
	native_reconfig_writedata_27,
	native_reconfig_writedata_28,
	native_reconfig_writedata_29,
	native_reconfig_writedata_30,
	native_reconfig_writedata_31,
	native_reconfig_write_1,
	native_reconfig_read_1,
	native_reconfig_address_12,
	native_reconfig_address_13,
	native_reconfig_address_14,
	native_reconfig_address_15,
	native_reconfig_address_16,
	native_reconfig_address_17,
	native_reconfig_address_18,
	native_reconfig_address_19,
	native_reconfig_address_20,
	native_reconfig_address_21,
	native_reconfig_address_22,
	native_reconfig_address_23,
	pif_testbus_sel_12,
	pif_testbus_sel_13,
	pif_testbus_sel_14,
	pif_testbus_sel_15,
	mutex_grant3,
	mutex_grant4,
	lif_waitrequest1,
	master_read,
	wbasic_read_82,
	lif_waitrequest2,
	basic_reconfig_waitrequest2,
	wbasic_writedata_1_8,
	wbasic_writedata_2_8,
	wbasic_writedata_0_8,
	wbasic_writedata_3_8,
	wbasic_writedata_4_8,
	wbasic_writedata_5_8,
	wbasic_writedata_6_8,
	wbasic_writedata_7_8,
	wbasic_writedata_8_8,
	wbasic_writedata_9_8,
	wbasic_writedata_10_8,
	wbasic_writedata_11_8,
	master_writedata_121,
	master_write_data_12,
	master_writedata_122,
	master_writedata_131,
	master_write_data_13,
	master_writedata_132,
	master_writedata_141,
	master_write_data_14,
	master_writedata_142,
	master_writedata_151,
	master_write_data_15,
	master_writedata_152,
	LessThan0,
	wbasic_write_83,
	lif_is_active,
	out_narrow_0,
	out_narrow_1,
	out_narrow_2,
	out_narrow_3,
	GND_port,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_16,
	reconfig_from_xcvr_0,
	reconfig_from_xcvr_46,
	reconfig_mgmt_writedata_17,
	reconfig_from_xcvr_1,
	reconfig_from_xcvr_47,
	reconfig_mgmt_writedata_18,
	reconfig_from_xcvr_2,
	reconfig_from_xcvr_48,
	reconfig_mgmt_writedata_19,
	reconfig_from_xcvr_3,
	reconfig_from_xcvr_49,
	reconfig_mgmt_writedata_20,
	reconfig_from_xcvr_4,
	reconfig_from_xcvr_50,
	reconfig_mgmt_writedata_21,
	reconfig_from_xcvr_5,
	reconfig_from_xcvr_51,
	reconfig_mgmt_writedata_22,
	reconfig_from_xcvr_6,
	reconfig_from_xcvr_52,
	reconfig_mgmt_writedata_23,
	reconfig_from_xcvr_7,
	reconfig_from_xcvr_53,
	reconfig_mgmt_writedata_24,
	reconfig_from_xcvr_8,
	reconfig_from_xcvr_54,
	reconfig_mgmt_writedata_25,
	reconfig_from_xcvr_9,
	reconfig_from_xcvr_55,
	reconfig_mgmt_writedata_26,
	reconfig_from_xcvr_10,
	reconfig_from_xcvr_56,
	reconfig_mgmt_writedata_27,
	reconfig_from_xcvr_11,
	reconfig_from_xcvr_57,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_from_xcvr_12,
	reconfig_from_xcvr_58,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_from_xcvr_13,
	reconfig_from_xcvr_59,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_from_xcvr_14,
	reconfig_from_xcvr_60,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15,
	reconfig_from_xcvr_15,
	reconfig_from_xcvr_61,
	reconfig_from_xcvr_24,
	reconfig_from_xcvr_70,
	reconfig_from_xcvr_16,
	reconfig_from_xcvr_62,
	reconfig_from_xcvr_32,
	reconfig_from_xcvr_78,
	reconfig_from_xcvr_25,
	reconfig_from_xcvr_71,
	reconfig_from_xcvr_17,
	reconfig_from_xcvr_63,
	reconfig_from_xcvr_33,
	reconfig_from_xcvr_79,
	reconfig_from_xcvr_26,
	reconfig_from_xcvr_72,
	reconfig_from_xcvr_18,
	reconfig_from_xcvr_64,
	reconfig_from_xcvr_34,
	reconfig_from_xcvr_80,
	reconfig_from_xcvr_27,
	reconfig_from_xcvr_73,
	reconfig_from_xcvr_19,
	reconfig_from_xcvr_65,
	reconfig_from_xcvr_35,
	reconfig_from_xcvr_81)/* synthesis synthesis_greybox=0 */;
output 	basic_reconfig_readdata_12;
output 	basic_reconfig_readdata_13;
output 	basic_reconfig_readdata_14;
output 	basic_reconfig_readdata_15;
output 	basic_reconfig_readdata_16;
output 	basic_reconfig_readdata_17;
output 	basic_reconfig_readdata_18;
output 	basic_reconfig_readdata_19;
output 	basic_reconfig_readdata_20;
output 	basic_reconfig_readdata_21;
output 	basic_reconfig_readdata_22;
output 	basic_reconfig_readdata_23;
output 	basic_reconfig_readdata_24;
output 	basic_reconfig_readdata_25;
output 	basic_reconfig_readdata_26;
output 	basic_reconfig_readdata_27;
output 	basic_reconfig_readdata_28;
output 	basic_reconfig_readdata_29;
output 	basic_reconfig_readdata_30;
output 	basic_reconfig_readdata_31;
input 	master_writedata_16;
input 	master_writedata_17;
input 	master_writedata_18;
input 	master_writedata_19;
input 	master_writedata_20;
input 	master_writedata_21;
input 	master_writedata_22;
input 	master_writedata_23;
input 	master_writedata_24;
input 	master_writedata_25;
input 	master_writedata_26;
input 	master_writedata_27;
input 	master_writedata_28;
input 	master_writedata_12;
input 	master_writedata_29;
input 	master_writedata_13;
input 	master_writedata_30;
input 	master_writedata_14;
input 	master_writedata_31;
input 	master_writedata_15;
output 	basic_reconfig_readdata_0;
output 	basic_reconfig_readdata_1;
output 	basic_reconfig_readdata_2;
output 	basic_reconfig_readdata_3;
output 	basic_reconfig_readdata_4;
output 	basic_reconfig_readdata_5;
input 	Equal2;
output 	basic_reconfig_readdata_6;
output 	basic_reconfig_readdata_7;
output 	basic_reconfig_readdata_8;
output 	basic_reconfig_readdata_9;
output 	basic_reconfig_readdata_10;
output 	basic_reconfig_readdata_11;
input 	mutex_grant;
input 	master_write;
input 	wbasic_write_8;
input 	wbasic_write_81;
input 	wbasic_write_82;
input 	mutex_grant1;
input 	wbasic_address_2_8;
input 	mutex_grant2;
input 	wbasic_address_0_8;
input 	wbasic_address_1_8;
output 	lif_waitrequest;
input 	wbasic_read_8;
input 	wbasic_read_81;
output 	basic_reconfig_waitrequest;
output 	basic_reconfig_waitrequest1;
input 	resync_chains0sync_r_1;
output 	native_reconfig_writedata_0;
output 	native_reconfig_writedata_1;
output 	native_reconfig_writedata_2;
output 	native_reconfig_writedata_3;
output 	native_reconfig_writedata_4;
output 	native_reconfig_writedata_5;
output 	native_reconfig_writedata_6;
output 	native_reconfig_writedata_7;
output 	native_reconfig_writedata_8;
output 	native_reconfig_writedata_9;
output 	native_reconfig_writedata_10;
output 	native_reconfig_writedata_11;
output 	native_reconfig_writedata_12;
output 	native_reconfig_writedata_13;
output 	native_reconfig_writedata_14;
output 	native_reconfig_writedata_15;
output 	native_reconfig_write_0;
output 	native_reconfig_read_0;
output 	native_reconfig_address_0;
output 	native_reconfig_address_1;
output 	native_reconfig_address_2;
output 	native_reconfig_address_3;
output 	native_reconfig_address_4;
output 	native_reconfig_address_5;
output 	native_reconfig_address_6;
output 	native_reconfig_address_7;
output 	native_reconfig_address_8;
output 	native_reconfig_address_9;
output 	native_reconfig_address_10;
output 	native_reconfig_address_11;
output 	pif_testbus_sel_0;
output 	pif_testbus_sel_1;
output 	pif_testbus_sel_2;
output 	pif_testbus_sel_3;
output 	pif_interface_sel;
output 	pif_ser_shift_load;
output 	native_reconfig_writedata_16;
output 	native_reconfig_writedata_17;
output 	native_reconfig_writedata_18;
output 	native_reconfig_writedata_19;
output 	native_reconfig_writedata_20;
output 	native_reconfig_writedata_21;
output 	native_reconfig_writedata_22;
output 	native_reconfig_writedata_23;
output 	native_reconfig_writedata_24;
output 	native_reconfig_writedata_25;
output 	native_reconfig_writedata_26;
output 	native_reconfig_writedata_27;
output 	native_reconfig_writedata_28;
output 	native_reconfig_writedata_29;
output 	native_reconfig_writedata_30;
output 	native_reconfig_writedata_31;
output 	native_reconfig_write_1;
output 	native_reconfig_read_1;
output 	native_reconfig_address_12;
output 	native_reconfig_address_13;
output 	native_reconfig_address_14;
output 	native_reconfig_address_15;
output 	native_reconfig_address_16;
output 	native_reconfig_address_17;
output 	native_reconfig_address_18;
output 	native_reconfig_address_19;
output 	native_reconfig_address_20;
output 	native_reconfig_address_21;
output 	native_reconfig_address_22;
output 	native_reconfig_address_23;
output 	pif_testbus_sel_12;
output 	pif_testbus_sel_13;
output 	pif_testbus_sel_14;
output 	pif_testbus_sel_15;
input 	mutex_grant3;
input 	mutex_grant4;
output 	lif_waitrequest1;
input 	master_read;
input 	wbasic_read_82;
output 	lif_waitrequest2;
output 	basic_reconfig_waitrequest2;
input 	wbasic_writedata_1_8;
input 	wbasic_writedata_2_8;
input 	wbasic_writedata_0_8;
input 	wbasic_writedata_3_8;
input 	wbasic_writedata_4_8;
input 	wbasic_writedata_5_8;
input 	wbasic_writedata_6_8;
input 	wbasic_writedata_7_8;
input 	wbasic_writedata_8_8;
input 	wbasic_writedata_9_8;
input 	wbasic_writedata_10_8;
input 	wbasic_writedata_11_8;
input 	master_writedata_121;
input 	master_write_data_12;
input 	master_writedata_122;
input 	master_writedata_131;
input 	master_write_data_13;
input 	master_writedata_132;
input 	master_writedata_141;
input 	master_write_data_14;
input 	master_writedata_142;
input 	master_writedata_151;
input 	master_write_data_15;
input 	master_writedata_152;
output 	LessThan0;
input 	wbasic_write_83;
input 	lif_is_active;
output 	out_narrow_0;
output 	out_narrow_1;
output 	out_narrow_2;
output 	out_narrow_3;
input 	GND_port;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_from_xcvr_0;
input 	reconfig_from_xcvr_46;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_from_xcvr_1;
input 	reconfig_from_xcvr_47;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_from_xcvr_2;
input 	reconfig_from_xcvr_48;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_from_xcvr_3;
input 	reconfig_from_xcvr_49;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_from_xcvr_4;
input 	reconfig_from_xcvr_50;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_from_xcvr_5;
input 	reconfig_from_xcvr_51;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_from_xcvr_6;
input 	reconfig_from_xcvr_52;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_from_xcvr_7;
input 	reconfig_from_xcvr_53;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_from_xcvr_8;
input 	reconfig_from_xcvr_54;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_from_xcvr_9;
input 	reconfig_from_xcvr_55;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_from_xcvr_10;
input 	reconfig_from_xcvr_56;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_from_xcvr_11;
input 	reconfig_from_xcvr_57;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_from_xcvr_12;
input 	reconfig_from_xcvr_58;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_from_xcvr_13;
input 	reconfig_from_xcvr_59;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_from_xcvr_14;
input 	reconfig_from_xcvr_60;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;
input 	reconfig_from_xcvr_15;
input 	reconfig_from_xcvr_61;
input 	reconfig_from_xcvr_24;
input 	reconfig_from_xcvr_70;
input 	reconfig_from_xcvr_16;
input 	reconfig_from_xcvr_62;
input 	reconfig_from_xcvr_32;
input 	reconfig_from_xcvr_78;
input 	reconfig_from_xcvr_25;
input 	reconfig_from_xcvr_71;
input 	reconfig_from_xcvr_17;
input 	reconfig_from_xcvr_63;
input 	reconfig_from_xcvr_33;
input 	reconfig_from_xcvr_79;
input 	reconfig_from_xcvr_26;
input 	reconfig_from_xcvr_72;
input 	reconfig_from_xcvr_18;
input 	reconfig_from_xcvr_64;
input 	reconfig_from_xcvr_34;
input 	reconfig_from_xcvr_80;
input 	reconfig_from_xcvr_27;
input 	reconfig_from_xcvr_73;
input 	reconfig_from_xcvr_19;
input 	reconfig_from_xcvr_65;
input 	reconfig_from_xcvr_35;
input 	reconfig_from_xcvr_81;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



RECONFIGURE_IP_av_xcvr_reconfig_basic a5(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.master_writedata_16(master_writedata_16),
	.master_writedata_17(master_writedata_17),
	.master_writedata_18(master_writedata_18),
	.master_writedata_19(master_writedata_19),
	.master_writedata_20(master_writedata_20),
	.master_writedata_21(master_writedata_21),
	.master_writedata_22(master_writedata_22),
	.master_writedata_23(master_writedata_23),
	.master_writedata_24(master_writedata_24),
	.master_writedata_25(master_writedata_25),
	.master_writedata_26(master_writedata_26),
	.master_writedata_27(master_writedata_27),
	.master_writedata_28(master_writedata_28),
	.master_writedata_12(master_writedata_12),
	.master_writedata_29(master_writedata_29),
	.master_writedata_13(master_writedata_13),
	.master_writedata_30(master_writedata_30),
	.master_writedata_14(master_writedata_14),
	.master_writedata_31(master_writedata_31),
	.master_writedata_15(master_writedata_15),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.Equal2(Equal2),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.mutex_grant(mutex_grant),
	.master_write(master_write),
	.wbasic_write_8(wbasic_write_8),
	.wbasic_write_81(wbasic_write_81),
	.wbasic_write_82(wbasic_write_82),
	.mutex_grant1(mutex_grant1),
	.wbasic_address_2_8(wbasic_address_2_8),
	.mutex_grant2(mutex_grant2),
	.wbasic_address_0_8(wbasic_address_0_8),
	.wbasic_address_1_8(wbasic_address_1_8),
	.lif_waitrequest(lif_waitrequest),
	.wbasic_read_8(wbasic_read_8),
	.wbasic_read_81(wbasic_read_81),
	.basic_reconfig_waitrequest({basic_reconfig_waitrequest}),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.native_reconfig_writedata_0(native_reconfig_writedata_0),
	.native_reconfig_writedata_1(native_reconfig_writedata_1),
	.native_reconfig_writedata_2(native_reconfig_writedata_2),
	.native_reconfig_writedata_3(native_reconfig_writedata_3),
	.native_reconfig_writedata_4(native_reconfig_writedata_4),
	.native_reconfig_writedata_5(native_reconfig_writedata_5),
	.native_reconfig_writedata_6(native_reconfig_writedata_6),
	.native_reconfig_writedata_7(native_reconfig_writedata_7),
	.native_reconfig_writedata_8(native_reconfig_writedata_8),
	.native_reconfig_writedata_9(native_reconfig_writedata_9),
	.native_reconfig_writedata_10(native_reconfig_writedata_10),
	.native_reconfig_writedata_11(native_reconfig_writedata_11),
	.native_reconfig_writedata_12(native_reconfig_writedata_12),
	.native_reconfig_writedata_13(native_reconfig_writedata_13),
	.native_reconfig_writedata_14(native_reconfig_writedata_14),
	.native_reconfig_writedata_15(native_reconfig_writedata_15),
	.native_reconfig_write_0(native_reconfig_write_0),
	.native_reconfig_read_0(native_reconfig_read_0),
	.native_reconfig_address_0(native_reconfig_address_0),
	.native_reconfig_address_1(native_reconfig_address_1),
	.native_reconfig_address_2(native_reconfig_address_2),
	.native_reconfig_address_3(native_reconfig_address_3),
	.native_reconfig_address_4(native_reconfig_address_4),
	.native_reconfig_address_5(native_reconfig_address_5),
	.native_reconfig_address_6(native_reconfig_address_6),
	.native_reconfig_address_7(native_reconfig_address_7),
	.native_reconfig_address_8(native_reconfig_address_8),
	.native_reconfig_address_9(native_reconfig_address_9),
	.native_reconfig_address_10(native_reconfig_address_10),
	.native_reconfig_address_11(native_reconfig_address_11),
	.pif_testbus_sel_0(pif_testbus_sel_0),
	.pif_testbus_sel_1(pif_testbus_sel_1),
	.pif_testbus_sel_2(pif_testbus_sel_2),
	.pif_testbus_sel_3(pif_testbus_sel_3),
	.pif_interface_sel1(pif_interface_sel),
	.pif_ser_shift_load1(pif_ser_shift_load),
	.native_reconfig_writedata_16(native_reconfig_writedata_16),
	.native_reconfig_writedata_17(native_reconfig_writedata_17),
	.native_reconfig_writedata_18(native_reconfig_writedata_18),
	.native_reconfig_writedata_19(native_reconfig_writedata_19),
	.native_reconfig_writedata_20(native_reconfig_writedata_20),
	.native_reconfig_writedata_21(native_reconfig_writedata_21),
	.native_reconfig_writedata_22(native_reconfig_writedata_22),
	.native_reconfig_writedata_23(native_reconfig_writedata_23),
	.native_reconfig_writedata_24(native_reconfig_writedata_24),
	.native_reconfig_writedata_25(native_reconfig_writedata_25),
	.native_reconfig_writedata_26(native_reconfig_writedata_26),
	.native_reconfig_writedata_27(native_reconfig_writedata_27),
	.native_reconfig_writedata_28(native_reconfig_writedata_28),
	.native_reconfig_writedata_29(native_reconfig_writedata_29),
	.native_reconfig_writedata_30(native_reconfig_writedata_30),
	.native_reconfig_writedata_31(native_reconfig_writedata_31),
	.native_reconfig_write_1(native_reconfig_write_1),
	.native_reconfig_read_1(native_reconfig_read_1),
	.native_reconfig_address_12(native_reconfig_address_12),
	.native_reconfig_address_13(native_reconfig_address_13),
	.native_reconfig_address_14(native_reconfig_address_14),
	.native_reconfig_address_15(native_reconfig_address_15),
	.native_reconfig_address_16(native_reconfig_address_16),
	.native_reconfig_address_17(native_reconfig_address_17),
	.native_reconfig_address_18(native_reconfig_address_18),
	.native_reconfig_address_19(native_reconfig_address_19),
	.native_reconfig_address_20(native_reconfig_address_20),
	.native_reconfig_address_21(native_reconfig_address_21),
	.native_reconfig_address_22(native_reconfig_address_22),
	.native_reconfig_address_23(native_reconfig_address_23),
	.pif_testbus_sel_12(pif_testbus_sel_12),
	.pif_testbus_sel_13(pif_testbus_sel_13),
	.pif_testbus_sel_14(pif_testbus_sel_14),
	.pif_testbus_sel_15(pif_testbus_sel_15),
	.mutex_grant3(mutex_grant3),
	.mutex_grant4(mutex_grant4),
	.lif_waitrequest1(lif_waitrequest1),
	.master_read(master_read),
	.wbasic_read_82(wbasic_read_82),
	.lif_waitrequest2(lif_waitrequest2),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.wbasic_writedata_1_8(wbasic_writedata_1_8),
	.wbasic_writedata_2_8(wbasic_writedata_2_8),
	.wbasic_writedata_0_8(wbasic_writedata_0_8),
	.wbasic_writedata_3_8(wbasic_writedata_3_8),
	.wbasic_writedata_4_8(wbasic_writedata_4_8),
	.wbasic_writedata_5_8(wbasic_writedata_5_8),
	.wbasic_writedata_6_8(wbasic_writedata_6_8),
	.wbasic_writedata_7_8(wbasic_writedata_7_8),
	.wbasic_writedata_8_8(wbasic_writedata_8_8),
	.wbasic_writedata_9_8(wbasic_writedata_9_8),
	.wbasic_writedata_10_8(wbasic_writedata_10_8),
	.wbasic_writedata_11_8(wbasic_writedata_11_8),
	.master_writedata_121(master_writedata_121),
	.master_write_data_12(master_write_data_12),
	.master_writedata_122(master_writedata_122),
	.master_writedata_131(master_writedata_131),
	.master_write_data_13(master_write_data_13),
	.master_writedata_132(master_writedata_132),
	.master_writedata_141(master_writedata_141),
	.master_write_data_14(master_write_data_14),
	.master_writedata_142(master_writedata_142),
	.master_writedata_151(master_writedata_151),
	.master_write_data_15(master_write_data_15),
	.master_writedata_152(master_writedata_152),
	.LessThan0(LessThan0),
	.wbasic_write_83(wbasic_write_83),
	.lif_is_active(lif_is_active),
	.out_narrow_0(out_narrow_0),
	.out_narrow_1(out_narrow_1),
	.out_narrow_2(out_narrow_2),
	.out_narrow_3(out_narrow_3),
	.GND_port(GND_port),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_from_xcvr_0(reconfig_from_xcvr_0),
	.reconfig_from_xcvr_46(reconfig_from_xcvr_46),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_from_xcvr_1(reconfig_from_xcvr_1),
	.reconfig_from_xcvr_47(reconfig_from_xcvr_47),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_from_xcvr_2(reconfig_from_xcvr_2),
	.reconfig_from_xcvr_48(reconfig_from_xcvr_48),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_from_xcvr_3(reconfig_from_xcvr_3),
	.reconfig_from_xcvr_49(reconfig_from_xcvr_49),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_from_xcvr_4(reconfig_from_xcvr_4),
	.reconfig_from_xcvr_50(reconfig_from_xcvr_50),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_from_xcvr_5(reconfig_from_xcvr_5),
	.reconfig_from_xcvr_51(reconfig_from_xcvr_51),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_from_xcvr_6(reconfig_from_xcvr_6),
	.reconfig_from_xcvr_52(reconfig_from_xcvr_52),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_from_xcvr_7(reconfig_from_xcvr_7),
	.reconfig_from_xcvr_53(reconfig_from_xcvr_53),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_from_xcvr_8(reconfig_from_xcvr_8),
	.reconfig_from_xcvr_54(reconfig_from_xcvr_54),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_from_xcvr_9(reconfig_from_xcvr_9),
	.reconfig_from_xcvr_55(reconfig_from_xcvr_55),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_from_xcvr_10(reconfig_from_xcvr_10),
	.reconfig_from_xcvr_56(reconfig_from_xcvr_56),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_from_xcvr_11(reconfig_from_xcvr_11),
	.reconfig_from_xcvr_57(reconfig_from_xcvr_57),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_from_xcvr_12(reconfig_from_xcvr_12),
	.reconfig_from_xcvr_58(reconfig_from_xcvr_58),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_from_xcvr_13(reconfig_from_xcvr_13),
	.reconfig_from_xcvr_59(reconfig_from_xcvr_59),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_from_xcvr_14(reconfig_from_xcvr_14),
	.reconfig_from_xcvr_60(reconfig_from_xcvr_60),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15),
	.reconfig_from_xcvr_15(reconfig_from_xcvr_15),
	.reconfig_from_xcvr_61(reconfig_from_xcvr_61),
	.reconfig_from_xcvr_24(reconfig_from_xcvr_24),
	.reconfig_from_xcvr_70(reconfig_from_xcvr_70),
	.reconfig_from_xcvr_16(reconfig_from_xcvr_16),
	.reconfig_from_xcvr_62(reconfig_from_xcvr_62),
	.reconfig_from_xcvr_32(reconfig_from_xcvr_32),
	.reconfig_from_xcvr_78(reconfig_from_xcvr_78),
	.reconfig_from_xcvr_25(reconfig_from_xcvr_25),
	.reconfig_from_xcvr_71(reconfig_from_xcvr_71),
	.reconfig_from_xcvr_17(reconfig_from_xcvr_17),
	.reconfig_from_xcvr_63(reconfig_from_xcvr_63),
	.reconfig_from_xcvr_33(reconfig_from_xcvr_33),
	.reconfig_from_xcvr_79(reconfig_from_xcvr_79),
	.reconfig_from_xcvr_26(reconfig_from_xcvr_26),
	.reconfig_from_xcvr_72(reconfig_from_xcvr_72),
	.reconfig_from_xcvr_18(reconfig_from_xcvr_18),
	.reconfig_from_xcvr_64(reconfig_from_xcvr_64),
	.reconfig_from_xcvr_34(reconfig_from_xcvr_34),
	.reconfig_from_xcvr_80(reconfig_from_xcvr_80),
	.reconfig_from_xcvr_27(reconfig_from_xcvr_27),
	.reconfig_from_xcvr_73(reconfig_from_xcvr_73),
	.reconfig_from_xcvr_19(reconfig_from_xcvr_19),
	.reconfig_from_xcvr_65(reconfig_from_xcvr_65),
	.reconfig_from_xcvr_35(reconfig_from_xcvr_35),
	.reconfig_from_xcvr_81(reconfig_from_xcvr_81));

endmodule

module RECONFIGURE_IP_av_xcvr_reconfig_basic (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	Equal2,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	mutex_grant,
	master_write,
	wbasic_write_8,
	wbasic_write_81,
	wbasic_write_82,
	mutex_grant1,
	wbasic_address_2_8,
	mutex_grant2,
	wbasic_address_0_8,
	wbasic_address_1_8,
	lif_waitrequest,
	wbasic_read_8,
	wbasic_read_81,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	resync_chains0sync_r_1,
	native_reconfig_writedata_0,
	native_reconfig_writedata_1,
	native_reconfig_writedata_2,
	native_reconfig_writedata_3,
	native_reconfig_writedata_4,
	native_reconfig_writedata_5,
	native_reconfig_writedata_6,
	native_reconfig_writedata_7,
	native_reconfig_writedata_8,
	native_reconfig_writedata_9,
	native_reconfig_writedata_10,
	native_reconfig_writedata_11,
	native_reconfig_writedata_12,
	native_reconfig_writedata_13,
	native_reconfig_writedata_14,
	native_reconfig_writedata_15,
	native_reconfig_write_0,
	native_reconfig_read_0,
	native_reconfig_address_0,
	native_reconfig_address_1,
	native_reconfig_address_2,
	native_reconfig_address_3,
	native_reconfig_address_4,
	native_reconfig_address_5,
	native_reconfig_address_6,
	native_reconfig_address_7,
	native_reconfig_address_8,
	native_reconfig_address_9,
	native_reconfig_address_10,
	native_reconfig_address_11,
	pif_testbus_sel_0,
	pif_testbus_sel_1,
	pif_testbus_sel_2,
	pif_testbus_sel_3,
	pif_interface_sel1,
	pif_ser_shift_load1,
	native_reconfig_writedata_16,
	native_reconfig_writedata_17,
	native_reconfig_writedata_18,
	native_reconfig_writedata_19,
	native_reconfig_writedata_20,
	native_reconfig_writedata_21,
	native_reconfig_writedata_22,
	native_reconfig_writedata_23,
	native_reconfig_writedata_24,
	native_reconfig_writedata_25,
	native_reconfig_writedata_26,
	native_reconfig_writedata_27,
	native_reconfig_writedata_28,
	native_reconfig_writedata_29,
	native_reconfig_writedata_30,
	native_reconfig_writedata_31,
	native_reconfig_write_1,
	native_reconfig_read_1,
	native_reconfig_address_12,
	native_reconfig_address_13,
	native_reconfig_address_14,
	native_reconfig_address_15,
	native_reconfig_address_16,
	native_reconfig_address_17,
	native_reconfig_address_18,
	native_reconfig_address_19,
	native_reconfig_address_20,
	native_reconfig_address_21,
	native_reconfig_address_22,
	native_reconfig_address_23,
	pif_testbus_sel_12,
	pif_testbus_sel_13,
	pif_testbus_sel_14,
	pif_testbus_sel_15,
	mutex_grant3,
	mutex_grant4,
	lif_waitrequest1,
	master_read,
	wbasic_read_82,
	lif_waitrequest2,
	basic_reconfig_waitrequest2,
	wbasic_writedata_1_8,
	wbasic_writedata_2_8,
	wbasic_writedata_0_8,
	wbasic_writedata_3_8,
	wbasic_writedata_4_8,
	wbasic_writedata_5_8,
	wbasic_writedata_6_8,
	wbasic_writedata_7_8,
	wbasic_writedata_8_8,
	wbasic_writedata_9_8,
	wbasic_writedata_10_8,
	wbasic_writedata_11_8,
	master_writedata_121,
	master_write_data_12,
	master_writedata_122,
	master_writedata_131,
	master_write_data_13,
	master_writedata_132,
	master_writedata_141,
	master_write_data_14,
	master_writedata_142,
	master_writedata_151,
	master_write_data_15,
	master_writedata_152,
	LessThan0,
	wbasic_write_83,
	lif_is_active,
	out_narrow_0,
	out_narrow_1,
	out_narrow_2,
	out_narrow_3,
	GND_port,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_16,
	reconfig_from_xcvr_0,
	reconfig_from_xcvr_46,
	reconfig_mgmt_writedata_17,
	reconfig_from_xcvr_1,
	reconfig_from_xcvr_47,
	reconfig_mgmt_writedata_18,
	reconfig_from_xcvr_2,
	reconfig_from_xcvr_48,
	reconfig_mgmt_writedata_19,
	reconfig_from_xcvr_3,
	reconfig_from_xcvr_49,
	reconfig_mgmt_writedata_20,
	reconfig_from_xcvr_4,
	reconfig_from_xcvr_50,
	reconfig_mgmt_writedata_21,
	reconfig_from_xcvr_5,
	reconfig_from_xcvr_51,
	reconfig_mgmt_writedata_22,
	reconfig_from_xcvr_6,
	reconfig_from_xcvr_52,
	reconfig_mgmt_writedata_23,
	reconfig_from_xcvr_7,
	reconfig_from_xcvr_53,
	reconfig_mgmt_writedata_24,
	reconfig_from_xcvr_8,
	reconfig_from_xcvr_54,
	reconfig_mgmt_writedata_25,
	reconfig_from_xcvr_9,
	reconfig_from_xcvr_55,
	reconfig_mgmt_writedata_26,
	reconfig_from_xcvr_10,
	reconfig_from_xcvr_56,
	reconfig_mgmt_writedata_27,
	reconfig_from_xcvr_11,
	reconfig_from_xcvr_57,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_from_xcvr_12,
	reconfig_from_xcvr_58,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_from_xcvr_13,
	reconfig_from_xcvr_59,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_from_xcvr_14,
	reconfig_from_xcvr_60,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15,
	reconfig_from_xcvr_15,
	reconfig_from_xcvr_61,
	reconfig_from_xcvr_24,
	reconfig_from_xcvr_70,
	reconfig_from_xcvr_16,
	reconfig_from_xcvr_62,
	reconfig_from_xcvr_32,
	reconfig_from_xcvr_78,
	reconfig_from_xcvr_25,
	reconfig_from_xcvr_71,
	reconfig_from_xcvr_17,
	reconfig_from_xcvr_63,
	reconfig_from_xcvr_33,
	reconfig_from_xcvr_79,
	reconfig_from_xcvr_26,
	reconfig_from_xcvr_72,
	reconfig_from_xcvr_18,
	reconfig_from_xcvr_64,
	reconfig_from_xcvr_34,
	reconfig_from_xcvr_80,
	reconfig_from_xcvr_27,
	reconfig_from_xcvr_73,
	reconfig_from_xcvr_19,
	reconfig_from_xcvr_65,
	reconfig_from_xcvr_35,
	reconfig_from_xcvr_81)/* synthesis synthesis_greybox=0 */;
output 	basic_reconfig_readdata_12;
output 	basic_reconfig_readdata_13;
output 	basic_reconfig_readdata_14;
output 	basic_reconfig_readdata_15;
output 	basic_reconfig_readdata_16;
output 	basic_reconfig_readdata_17;
output 	basic_reconfig_readdata_18;
output 	basic_reconfig_readdata_19;
output 	basic_reconfig_readdata_20;
output 	basic_reconfig_readdata_21;
output 	basic_reconfig_readdata_22;
output 	basic_reconfig_readdata_23;
output 	basic_reconfig_readdata_24;
output 	basic_reconfig_readdata_25;
output 	basic_reconfig_readdata_26;
output 	basic_reconfig_readdata_27;
output 	basic_reconfig_readdata_28;
output 	basic_reconfig_readdata_29;
output 	basic_reconfig_readdata_30;
output 	basic_reconfig_readdata_31;
input 	master_writedata_16;
input 	master_writedata_17;
input 	master_writedata_18;
input 	master_writedata_19;
input 	master_writedata_20;
input 	master_writedata_21;
input 	master_writedata_22;
input 	master_writedata_23;
input 	master_writedata_24;
input 	master_writedata_25;
input 	master_writedata_26;
input 	master_writedata_27;
input 	master_writedata_28;
input 	master_writedata_12;
input 	master_writedata_29;
input 	master_writedata_13;
input 	master_writedata_30;
input 	master_writedata_14;
input 	master_writedata_31;
input 	master_writedata_15;
output 	basic_reconfig_readdata_0;
output 	basic_reconfig_readdata_1;
output 	basic_reconfig_readdata_2;
output 	basic_reconfig_readdata_3;
output 	basic_reconfig_readdata_4;
output 	basic_reconfig_readdata_5;
input 	Equal2;
output 	basic_reconfig_readdata_6;
output 	basic_reconfig_readdata_7;
output 	basic_reconfig_readdata_8;
output 	basic_reconfig_readdata_9;
output 	basic_reconfig_readdata_10;
output 	basic_reconfig_readdata_11;
input 	mutex_grant;
input 	master_write;
input 	wbasic_write_8;
input 	wbasic_write_81;
input 	wbasic_write_82;
input 	mutex_grant1;
input 	wbasic_address_2_8;
input 	mutex_grant2;
input 	wbasic_address_0_8;
input 	wbasic_address_1_8;
output 	lif_waitrequest;
input 	wbasic_read_8;
input 	wbasic_read_81;
output 	[0:0] basic_reconfig_waitrequest;
output 	basic_reconfig_waitrequest1;
input 	resync_chains0sync_r_1;
output 	native_reconfig_writedata_0;
output 	native_reconfig_writedata_1;
output 	native_reconfig_writedata_2;
output 	native_reconfig_writedata_3;
output 	native_reconfig_writedata_4;
output 	native_reconfig_writedata_5;
output 	native_reconfig_writedata_6;
output 	native_reconfig_writedata_7;
output 	native_reconfig_writedata_8;
output 	native_reconfig_writedata_9;
output 	native_reconfig_writedata_10;
output 	native_reconfig_writedata_11;
output 	native_reconfig_writedata_12;
output 	native_reconfig_writedata_13;
output 	native_reconfig_writedata_14;
output 	native_reconfig_writedata_15;
output 	native_reconfig_write_0;
output 	native_reconfig_read_0;
output 	native_reconfig_address_0;
output 	native_reconfig_address_1;
output 	native_reconfig_address_2;
output 	native_reconfig_address_3;
output 	native_reconfig_address_4;
output 	native_reconfig_address_5;
output 	native_reconfig_address_6;
output 	native_reconfig_address_7;
output 	native_reconfig_address_8;
output 	native_reconfig_address_9;
output 	native_reconfig_address_10;
output 	native_reconfig_address_11;
output 	pif_testbus_sel_0;
output 	pif_testbus_sel_1;
output 	pif_testbus_sel_2;
output 	pif_testbus_sel_3;
output 	pif_interface_sel1;
output 	pif_ser_shift_load1;
output 	native_reconfig_writedata_16;
output 	native_reconfig_writedata_17;
output 	native_reconfig_writedata_18;
output 	native_reconfig_writedata_19;
output 	native_reconfig_writedata_20;
output 	native_reconfig_writedata_21;
output 	native_reconfig_writedata_22;
output 	native_reconfig_writedata_23;
output 	native_reconfig_writedata_24;
output 	native_reconfig_writedata_25;
output 	native_reconfig_writedata_26;
output 	native_reconfig_writedata_27;
output 	native_reconfig_writedata_28;
output 	native_reconfig_writedata_29;
output 	native_reconfig_writedata_30;
output 	native_reconfig_writedata_31;
output 	native_reconfig_write_1;
output 	native_reconfig_read_1;
output 	native_reconfig_address_12;
output 	native_reconfig_address_13;
output 	native_reconfig_address_14;
output 	native_reconfig_address_15;
output 	native_reconfig_address_16;
output 	native_reconfig_address_17;
output 	native_reconfig_address_18;
output 	native_reconfig_address_19;
output 	native_reconfig_address_20;
output 	native_reconfig_address_21;
output 	native_reconfig_address_22;
output 	native_reconfig_address_23;
output 	pif_testbus_sel_12;
output 	pif_testbus_sel_13;
output 	pif_testbus_sel_14;
output 	pif_testbus_sel_15;
input 	mutex_grant3;
input 	mutex_grant4;
output 	lif_waitrequest1;
input 	master_read;
input 	wbasic_read_82;
output 	lif_waitrequest2;
output 	basic_reconfig_waitrequest2;
input 	wbasic_writedata_1_8;
input 	wbasic_writedata_2_8;
input 	wbasic_writedata_0_8;
input 	wbasic_writedata_3_8;
input 	wbasic_writedata_4_8;
input 	wbasic_writedata_5_8;
input 	wbasic_writedata_6_8;
input 	wbasic_writedata_7_8;
input 	wbasic_writedata_8_8;
input 	wbasic_writedata_9_8;
input 	wbasic_writedata_10_8;
input 	wbasic_writedata_11_8;
input 	master_writedata_121;
input 	master_write_data_12;
input 	master_writedata_122;
input 	master_writedata_131;
input 	master_write_data_13;
input 	master_writedata_132;
input 	master_writedata_141;
input 	master_write_data_14;
input 	master_writedata_142;
input 	master_writedata_151;
input 	master_write_data_15;
input 	master_writedata_152;
output 	LessThan0;
input 	wbasic_write_83;
input 	lif_is_active;
output 	out_narrow_0;
output 	out_narrow_1;
output 	out_narrow_2;
output 	out_narrow_3;
input 	GND_port;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_from_xcvr_0;
input 	reconfig_from_xcvr_46;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_from_xcvr_1;
input 	reconfig_from_xcvr_47;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_from_xcvr_2;
input 	reconfig_from_xcvr_48;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_from_xcvr_3;
input 	reconfig_from_xcvr_49;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_from_xcvr_4;
input 	reconfig_from_xcvr_50;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_from_xcvr_5;
input 	reconfig_from_xcvr_51;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_from_xcvr_6;
input 	reconfig_from_xcvr_52;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_from_xcvr_7;
input 	reconfig_from_xcvr_53;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_from_xcvr_8;
input 	reconfig_from_xcvr_54;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_from_xcvr_9;
input 	reconfig_from_xcvr_55;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_from_xcvr_10;
input 	reconfig_from_xcvr_56;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_from_xcvr_11;
input 	reconfig_from_xcvr_57;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_from_xcvr_12;
input 	reconfig_from_xcvr_58;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_from_xcvr_13;
input 	reconfig_from_xcvr_59;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_from_xcvr_14;
input 	reconfig_from_xcvr_60;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;
input 	reconfig_from_xcvr_15;
input 	reconfig_from_xcvr_61;
input 	reconfig_from_xcvr_24;
input 	reconfig_from_xcvr_70;
input 	reconfig_from_xcvr_16;
input 	reconfig_from_xcvr_62;
input 	reconfig_from_xcvr_32;
input 	reconfig_from_xcvr_78;
input 	reconfig_from_xcvr_25;
input 	reconfig_from_xcvr_71;
input 	reconfig_from_xcvr_17;
input 	reconfig_from_xcvr_63;
input 	reconfig_from_xcvr_33;
input 	reconfig_from_xcvr_79;
input 	reconfig_from_xcvr_26;
input 	reconfig_from_xcvr_72;
input 	reconfig_from_xcvr_18;
input 	reconfig_from_xcvr_64;
input 	reconfig_from_xcvr_34;
input 	reconfig_from_xcvr_80;
input 	reconfig_from_xcvr_27;
input 	reconfig_from_xcvr_73;
input 	reconfig_from_xcvr_19;
input 	reconfig_from_xcvr_65;
input 	reconfig_from_xcvr_35;
input 	reconfig_from_xcvr_81;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lif[0].logical_if|pif_ena[0]~q ;
wire \pif[0].pif_arb|grant[0]~q ;
wire \lif[0].logical_if|pif_ena[1]~q ;
wire \pif[1].pif_arb|grant[0]~q ;
wire \lif[0].logical_if|lif_csr|reg_plock~q ;
wire \Add0~41_sumout ;
wire \reg_init[9]~0_combout ;
wire \init_done~0_combout ;
wire \init_done~q ;
wire \always0~0_combout ;
wire \reg_init[0]~q ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \reg_init[1]~q ;
wire \Add0~46 ;
wire \Add0~37_sumout ;
wire \reg_init[2]~q ;
wire \Add0~38 ;
wire \Add0~25_sumout ;
wire \reg_init[3]~q ;
wire \Add0~26 ;
wire \Add0~33_sumout ;
wire \reg_init[4]~q ;
wire \Add0~34 ;
wire \Add0~29_sumout ;
wire \reg_init[5]~q ;
wire \Add0~30 ;
wire \Add0~5_sumout ;
wire \reg_init[6]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \reg_init[7]~q ;
wire \Add0~10 ;
wire \Add0~17_sumout ;
wire \reg_init[8]~q ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \reg_init[9]~q ;
wire \Add0~14 ;
wire \Add0~21_sumout ;
wire \reg_init[10]~q ;
wire \Add0~22 ;
wire \Add0~1_sumout ;
wire \reg_init[11]~q ;
wire \pif_ser_shift_load~0_combout ;
wire \pif_ser_shift_load~1_combout ;
wire \pif_ser_shift_load~2_combout ;


RECONFIGURE_IP_alt_xcvr_arbiter_2 \pif[1].pif_arb (
	.pif_ena_1(\lif[0].logical_if|pif_ena[1]~q ),
	.grant_0(\pif[1].pif_arb|grant[0]~q ),
	.reg_plock(\lif[0].logical_if|lif_csr|reg_plock~q ),
	.mgmt_clk_clk(mgmt_clk_clk));

RECONFIGURE_IP_alt_xcvr_arbiter_1 \pif[0].pif_arb (
	.pif_ena_0(\lif[0].logical_if|pif_ena[0]~q ),
	.grant_0(\pif[0].pif_arb|grant[0]~q ),
	.reg_plock(\lif[0].logical_if|lif_csr|reg_plock~q ),
	.mgmt_clk_clk(mgmt_clk_clk));

RECONFIGURE_IP_av_xrbasic_lif \lif[0].logical_if (
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.master_writedata_16(master_writedata_16),
	.master_writedata_17(master_writedata_17),
	.master_writedata_18(master_writedata_18),
	.master_writedata_19(master_writedata_19),
	.master_writedata_20(master_writedata_20),
	.master_writedata_21(master_writedata_21),
	.master_writedata_22(master_writedata_22),
	.master_writedata_23(master_writedata_23),
	.master_writedata_24(master_writedata_24),
	.master_writedata_25(master_writedata_25),
	.master_writedata_26(master_writedata_26),
	.master_writedata_27(master_writedata_27),
	.master_writedata_28(master_writedata_28),
	.master_writedata_12(master_writedata_12),
	.master_writedata_29(master_writedata_29),
	.master_writedata_13(master_writedata_13),
	.master_writedata_30(master_writedata_30),
	.master_writedata_14(master_writedata_14),
	.master_writedata_31(master_writedata_31),
	.master_writedata_15(master_writedata_15),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.Equal2(Equal2),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.mutex_grant(mutex_grant),
	.master_write(master_write),
	.wbasic_write_8(wbasic_write_8),
	.wbasic_write_81(wbasic_write_81),
	.wbasic_write_82(wbasic_write_82),
	.mutex_grant1(mutex_grant1),
	.wbasic_address_2_8(wbasic_address_2_8),
	.mutex_grant2(mutex_grant2),
	.wbasic_address_0_8(wbasic_address_0_8),
	.wbasic_address_1_8(wbasic_address_1_8),
	.lif_waitrequest(lif_waitrequest),
	.wbasic_read_8(wbasic_read_8),
	.wbasic_read_81(wbasic_read_81),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest[0]),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.pif_ena_0(\lif[0].logical_if|pif_ena[0]~q ),
	.grant_0(\pif[0].pif_arb|grant[0]~q ),
	.native_reconfig_writedata_0(native_reconfig_writedata_0),
	.native_reconfig_writedata_1(native_reconfig_writedata_1),
	.native_reconfig_writedata_2(native_reconfig_writedata_2),
	.native_reconfig_writedata_3(native_reconfig_writedata_3),
	.native_reconfig_writedata_4(native_reconfig_writedata_4),
	.native_reconfig_writedata_5(native_reconfig_writedata_5),
	.native_reconfig_writedata_6(native_reconfig_writedata_6),
	.native_reconfig_writedata_7(native_reconfig_writedata_7),
	.native_reconfig_writedata_8(native_reconfig_writedata_8),
	.native_reconfig_writedata_9(native_reconfig_writedata_9),
	.native_reconfig_writedata_10(native_reconfig_writedata_10),
	.native_reconfig_writedata_11(native_reconfig_writedata_11),
	.native_reconfig_writedata_12(native_reconfig_writedata_12),
	.native_reconfig_writedata_13(native_reconfig_writedata_13),
	.native_reconfig_writedata_14(native_reconfig_writedata_14),
	.native_reconfig_writedata_15(native_reconfig_writedata_15),
	.native_reconfig_write_0(native_reconfig_write_0),
	.native_reconfig_read_0(native_reconfig_read_0),
	.native_reconfig_address_0(native_reconfig_address_0),
	.native_reconfig_address_1(native_reconfig_address_1),
	.native_reconfig_address_2(native_reconfig_address_2),
	.native_reconfig_address_3(native_reconfig_address_3),
	.native_reconfig_address_4(native_reconfig_address_4),
	.native_reconfig_address_5(native_reconfig_address_5),
	.native_reconfig_address_6(native_reconfig_address_6),
	.native_reconfig_address_7(native_reconfig_address_7),
	.native_reconfig_address_8(native_reconfig_address_8),
	.native_reconfig_address_9(native_reconfig_address_9),
	.native_reconfig_address_10(native_reconfig_address_10),
	.native_reconfig_address_11(native_reconfig_address_11),
	.pif_testbus_sel_0(pif_testbus_sel_0),
	.pif_testbus_sel_1(pif_testbus_sel_1),
	.pif_testbus_sel_2(pif_testbus_sel_2),
	.pif_testbus_sel_3(pif_testbus_sel_3),
	.pif_ena_1(\lif[0].logical_if|pif_ena[1]~q ),
	.grant_01(\pif[1].pif_arb|grant[0]~q ),
	.native_reconfig_writedata_16(native_reconfig_writedata_16),
	.native_reconfig_writedata_17(native_reconfig_writedata_17),
	.native_reconfig_writedata_18(native_reconfig_writedata_18),
	.native_reconfig_writedata_19(native_reconfig_writedata_19),
	.native_reconfig_writedata_20(native_reconfig_writedata_20),
	.native_reconfig_writedata_21(native_reconfig_writedata_21),
	.native_reconfig_writedata_22(native_reconfig_writedata_22),
	.native_reconfig_writedata_23(native_reconfig_writedata_23),
	.native_reconfig_writedata_24(native_reconfig_writedata_24),
	.native_reconfig_writedata_25(native_reconfig_writedata_25),
	.native_reconfig_writedata_26(native_reconfig_writedata_26),
	.native_reconfig_writedata_27(native_reconfig_writedata_27),
	.native_reconfig_writedata_28(native_reconfig_writedata_28),
	.native_reconfig_writedata_29(native_reconfig_writedata_29),
	.native_reconfig_writedata_30(native_reconfig_writedata_30),
	.native_reconfig_writedata_31(native_reconfig_writedata_31),
	.native_reconfig_write_1(native_reconfig_write_1),
	.native_reconfig_read_1(native_reconfig_read_1),
	.native_reconfig_address_12(native_reconfig_address_12),
	.native_reconfig_address_13(native_reconfig_address_13),
	.native_reconfig_address_14(native_reconfig_address_14),
	.native_reconfig_address_15(native_reconfig_address_15),
	.native_reconfig_address_16(native_reconfig_address_16),
	.native_reconfig_address_17(native_reconfig_address_17),
	.native_reconfig_address_18(native_reconfig_address_18),
	.native_reconfig_address_19(native_reconfig_address_19),
	.native_reconfig_address_20(native_reconfig_address_20),
	.native_reconfig_address_21(native_reconfig_address_21),
	.native_reconfig_address_22(native_reconfig_address_22),
	.native_reconfig_address_23(native_reconfig_address_23),
	.pif_testbus_sel_12(pif_testbus_sel_12),
	.pif_testbus_sel_13(pif_testbus_sel_13),
	.pif_testbus_sel_14(pif_testbus_sel_14),
	.pif_testbus_sel_15(pif_testbus_sel_15),
	.reg_plock(\lif[0].logical_if|lif_csr|reg_plock~q ),
	.mutex_grant3(mutex_grant3),
	.mutex_grant4(mutex_grant4),
	.lif_waitrequest1(lif_waitrequest1),
	.master_read(master_read),
	.wbasic_read_82(wbasic_read_82),
	.lif_waitrequest2(lif_waitrequest2),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.wbasic_writedata_1_8(wbasic_writedata_1_8),
	.wbasic_writedata_2_8(wbasic_writedata_2_8),
	.wbasic_writedata_0_8(wbasic_writedata_0_8),
	.wbasic_writedata_3_8(wbasic_writedata_3_8),
	.wbasic_writedata_4_8(wbasic_writedata_4_8),
	.wbasic_writedata_5_8(wbasic_writedata_5_8),
	.wbasic_writedata_6_8(wbasic_writedata_6_8),
	.wbasic_writedata_7_8(wbasic_writedata_7_8),
	.wbasic_writedata_8_8(wbasic_writedata_8_8),
	.wbasic_writedata_9_8(wbasic_writedata_9_8),
	.wbasic_writedata_10_8(wbasic_writedata_10_8),
	.wbasic_writedata_11_8(wbasic_writedata_11_8),
	.master_writedata_121(master_writedata_121),
	.master_write_data_12(master_write_data_12),
	.master_writedata_122(master_writedata_122),
	.master_writedata_131(master_writedata_131),
	.master_write_data_13(master_write_data_13),
	.master_writedata_132(master_writedata_132),
	.master_writedata_141(master_writedata_141),
	.master_write_data_14(master_write_data_14),
	.master_writedata_142(master_writedata_142),
	.master_writedata_151(master_writedata_151),
	.master_write_data_15(master_write_data_15),
	.master_writedata_152(master_writedata_152),
	.wbasic_write_83(wbasic_write_83),
	.lif_is_active(lif_is_active),
	.out_narrow_0(out_narrow_0),
	.out_narrow_1(out_narrow_1),
	.out_narrow_2(out_narrow_2),
	.out_narrow_3(out_narrow_3),
	.GND_port(GND_port),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_from_xcvr_0(reconfig_from_xcvr_0),
	.reconfig_from_xcvr_46(reconfig_from_xcvr_46),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_from_xcvr_1(reconfig_from_xcvr_1),
	.reconfig_from_xcvr_47(reconfig_from_xcvr_47),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_from_xcvr_2(reconfig_from_xcvr_2),
	.reconfig_from_xcvr_48(reconfig_from_xcvr_48),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_from_xcvr_3(reconfig_from_xcvr_3),
	.reconfig_from_xcvr_49(reconfig_from_xcvr_49),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_from_xcvr_4(reconfig_from_xcvr_4),
	.reconfig_from_xcvr_50(reconfig_from_xcvr_50),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_from_xcvr_5(reconfig_from_xcvr_5),
	.reconfig_from_xcvr_51(reconfig_from_xcvr_51),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_from_xcvr_6(reconfig_from_xcvr_6),
	.reconfig_from_xcvr_52(reconfig_from_xcvr_52),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_from_xcvr_7(reconfig_from_xcvr_7),
	.reconfig_from_xcvr_53(reconfig_from_xcvr_53),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_from_xcvr_8(reconfig_from_xcvr_8),
	.reconfig_from_xcvr_54(reconfig_from_xcvr_54),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_from_xcvr_9(reconfig_from_xcvr_9),
	.reconfig_from_xcvr_55(reconfig_from_xcvr_55),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_from_xcvr_10(reconfig_from_xcvr_10),
	.reconfig_from_xcvr_56(reconfig_from_xcvr_56),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_from_xcvr_11(reconfig_from_xcvr_11),
	.reconfig_from_xcvr_57(reconfig_from_xcvr_57),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_from_xcvr_12(reconfig_from_xcvr_12),
	.reconfig_from_xcvr_58(reconfig_from_xcvr_58),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_from_xcvr_13(reconfig_from_xcvr_13),
	.reconfig_from_xcvr_59(reconfig_from_xcvr_59),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_from_xcvr_14(reconfig_from_xcvr_14),
	.reconfig_from_xcvr_60(reconfig_from_xcvr_60),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15),
	.reconfig_from_xcvr_15(reconfig_from_xcvr_15),
	.reconfig_from_xcvr_61(reconfig_from_xcvr_61),
	.reconfig_from_xcvr_24(reconfig_from_xcvr_24),
	.reconfig_from_xcvr_70(reconfig_from_xcvr_70),
	.reconfig_from_xcvr_16(reconfig_from_xcvr_16),
	.reconfig_from_xcvr_62(reconfig_from_xcvr_62),
	.reconfig_from_xcvr_32(reconfig_from_xcvr_32),
	.reconfig_from_xcvr_78(reconfig_from_xcvr_78),
	.reconfig_from_xcvr_25(reconfig_from_xcvr_25),
	.reconfig_from_xcvr_71(reconfig_from_xcvr_71),
	.reconfig_from_xcvr_17(reconfig_from_xcvr_17),
	.reconfig_from_xcvr_63(reconfig_from_xcvr_63),
	.reconfig_from_xcvr_33(reconfig_from_xcvr_33),
	.reconfig_from_xcvr_79(reconfig_from_xcvr_79),
	.reconfig_from_xcvr_26(reconfig_from_xcvr_26),
	.reconfig_from_xcvr_72(reconfig_from_xcvr_72),
	.reconfig_from_xcvr_18(reconfig_from_xcvr_18),
	.reconfig_from_xcvr_64(reconfig_from_xcvr_64),
	.reconfig_from_xcvr_34(reconfig_from_xcvr_34),
	.reconfig_from_xcvr_80(reconfig_from_xcvr_80),
	.reconfig_from_xcvr_27(reconfig_from_xcvr_27),
	.reconfig_from_xcvr_73(reconfig_from_xcvr_73),
	.reconfig_from_xcvr_19(reconfig_from_xcvr_19),
	.reconfig_from_xcvr_65(reconfig_from_xcvr_65),
	.reconfig_from_xcvr_35(reconfig_from_xcvr_35),
	.reconfig_from_xcvr_81(reconfig_from_xcvr_81));

dffeas pif_interface_sel(
	.clk(mgmt_clk_clk),
	.d(LessThan0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pif_interface_sel1),
	.prn(vcc));
defparam pif_interface_sel.is_wysiwyg = "true";
defparam pif_interface_sel.power_up = "low";

dffeas pif_ser_shift_load(
	.clk(mgmt_clk_clk),
	.d(\pif_ser_shift_load~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pif_ser_shift_load1),
	.prn(vcc));
defparam pif_ser_shift_load.is_wysiwyg = "true";
defparam pif_ser_shift_load.power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\reg_init[11]~q ),
	.datab(!\reg_init[6]~q ),
	.datac(!\reg_init[7]~q ),
	.datad(!\reg_init[9]~q ),
	.datae(!\reg_init[8]~q ),
	.dataf(!\reg_init[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h0155555555555555;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \reg_init[9]~0 (
	.dataa(!LessThan0),
	.datab(!\always0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_init[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_init[9]~0 .extended_lut = "off";
defparam \reg_init[9]~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \reg_init[9]~0 .shared_arith = "off";

cyclonev_lcell_comb \init_done~0 (
	.dataa(!\init_done~q ),
	.datab(!\reg_init[9]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\init_done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \init_done~0 .extended_lut = "off";
defparam \init_done~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \init_done~0 .shared_arith = "off";

dffeas init_done(
	.clk(mgmt_clk_clk),
	.d(\init_done~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\init_done~q ),
	.prn(vcc));
defparam init_done.is_wysiwyg = "true";
defparam init_done.power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!resync_chains0sync_r_1),
	.datab(!\init_done~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8888888888888888;
defparam \always0~0 .shared_arith = "off";

dffeas \reg_init[0] (
	.clk(mgmt_clk_clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[0]~q ),
	.prn(vcc));
defparam \reg_init[0] .is_wysiwyg = "true";
defparam \reg_init[0] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \reg_init[1] (
	.clk(mgmt_clk_clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[1]~q ),
	.prn(vcc));
defparam \reg_init[1] .is_wysiwyg = "true";
defparam \reg_init[1] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \reg_init[2] (
	.clk(mgmt_clk_clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[2]~q ),
	.prn(vcc));
defparam \reg_init[2] .is_wysiwyg = "true";
defparam \reg_init[2] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \reg_init[3] (
	.clk(mgmt_clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[3]~q ),
	.prn(vcc));
defparam \reg_init[3] .is_wysiwyg = "true";
defparam \reg_init[3] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \reg_init[4] (
	.clk(mgmt_clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[4]~q ),
	.prn(vcc));
defparam \reg_init[4] .is_wysiwyg = "true";
defparam \reg_init[4] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \reg_init[5] (
	.clk(mgmt_clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[5]~q ),
	.prn(vcc));
defparam \reg_init[5] .is_wysiwyg = "true";
defparam \reg_init[5] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \reg_init[6] (
	.clk(mgmt_clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[6]~q ),
	.prn(vcc));
defparam \reg_init[6] .is_wysiwyg = "true";
defparam \reg_init[6] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \reg_init[7] (
	.clk(mgmt_clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[7]~q ),
	.prn(vcc));
defparam \reg_init[7] .is_wysiwyg = "true";
defparam \reg_init[7] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \reg_init[8] (
	.clk(mgmt_clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[8]~q ),
	.prn(vcc));
defparam \reg_init[8] .is_wysiwyg = "true";
defparam \reg_init[8] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \reg_init[9] (
	.clk(mgmt_clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[9]~q ),
	.prn(vcc));
defparam \reg_init[9] .is_wysiwyg = "true";
defparam \reg_init[9] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \reg_init[10] (
	.clk(mgmt_clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[10]~q ),
	.prn(vcc));
defparam \reg_init[10] .is_wysiwyg = "true";
defparam \reg_init[10] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_init[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \reg_init[11] (
	.clk(mgmt_clk_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\reg_init[9]~0_combout ),
	.q(\reg_init[11]~q ),
	.prn(vcc));
defparam \reg_init[11] .is_wysiwyg = "true";
defparam \reg_init[11] .power_up = "low";

cyclonev_lcell_comb \pif_ser_shift_load~0 (
	.dataa(!\reg_init[6]~q ),
	.datab(!\reg_init[7]~q ),
	.datac(!\reg_init[5]~q ),
	.datad(!\reg_init[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_ser_shift_load~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_ser_shift_load~0 .extended_lut = "off";
defparam \pif_ser_shift_load~0 .lut_mask = 64'h0002000200020002;
defparam \pif_ser_shift_load~0 .shared_arith = "off";

cyclonev_lcell_comb \pif_ser_shift_load~1 (
	.dataa(!\reg_init[9]~q ),
	.datab(!\reg_init[8]~q ),
	.datac(!\reg_init[10]~q ),
	.datad(!\reg_init[2]~q ),
	.datae(!\reg_init[0]~q ),
	.dataf(!\reg_init[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_ser_shift_load~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_ser_shift_load~1 .extended_lut = "off";
defparam \pif_ser_shift_load~1 .lut_mask = 64'h0080008000808000;
defparam \pif_ser_shift_load~1 .shared_arith = "off";

cyclonev_lcell_comb \pif_ser_shift_load~2 (
	.dataa(!\reg_init[11]~q ),
	.datab(!\reg_init[3]~q ),
	.datac(!\pif_ser_shift_load~0_combout ),
	.datad(!\pif_ser_shift_load~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_ser_shift_load~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_ser_shift_load~2 .extended_lut = "off";
defparam \pif_ser_shift_load~2 .lut_mask = 64'h0001000100010001;
defparam \pif_ser_shift_load~2 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_arbiter_1 (
	pif_ena_0,
	grant_0,
	reg_plock,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	pif_ena_0;
output 	grant_0;
input 	reg_plock;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \grant[0]~0_combout ;


dffeas \grant[0] (
	.clk(mgmt_clk_clk),
	.d(\grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(grant_0),
	.prn(vcc));
defparam \grant[0] .is_wysiwyg = "true";
defparam \grant[0] .power_up = "low";

cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!reg_plock),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'h3737373737373737;
defparam \grant[0]~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_arbiter_2 (
	pif_ena_1,
	grant_0,
	reg_plock,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	pif_ena_1;
output 	grant_0;
input 	reg_plock;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \grant[0]~0_combout ;


dffeas \grant[0] (
	.clk(mgmt_clk_clk),
	.d(\grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(grant_0),
	.prn(vcc));
defparam \grant[0] .is_wysiwyg = "true";
defparam \grant[0] .power_up = "low";

cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!pif_ena_1),
	.datab(!grant_0),
	.datac(!reg_plock),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\grant[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'h3737373737373737;
defparam \grant[0]~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_av_xrbasic_lif (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	Equal2,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	mutex_grant,
	master_write,
	wbasic_write_8,
	wbasic_write_81,
	wbasic_write_82,
	mutex_grant1,
	wbasic_address_2_8,
	mutex_grant2,
	wbasic_address_0_8,
	wbasic_address_1_8,
	lif_waitrequest,
	wbasic_read_8,
	wbasic_read_81,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	resync_chains0sync_r_1,
	pif_ena_0,
	grant_0,
	native_reconfig_writedata_0,
	native_reconfig_writedata_1,
	native_reconfig_writedata_2,
	native_reconfig_writedata_3,
	native_reconfig_writedata_4,
	native_reconfig_writedata_5,
	native_reconfig_writedata_6,
	native_reconfig_writedata_7,
	native_reconfig_writedata_8,
	native_reconfig_writedata_9,
	native_reconfig_writedata_10,
	native_reconfig_writedata_11,
	native_reconfig_writedata_12,
	native_reconfig_writedata_13,
	native_reconfig_writedata_14,
	native_reconfig_writedata_15,
	native_reconfig_write_0,
	native_reconfig_read_0,
	native_reconfig_address_0,
	native_reconfig_address_1,
	native_reconfig_address_2,
	native_reconfig_address_3,
	native_reconfig_address_4,
	native_reconfig_address_5,
	native_reconfig_address_6,
	native_reconfig_address_7,
	native_reconfig_address_8,
	native_reconfig_address_9,
	native_reconfig_address_10,
	native_reconfig_address_11,
	pif_testbus_sel_0,
	pif_testbus_sel_1,
	pif_testbus_sel_2,
	pif_testbus_sel_3,
	pif_ena_1,
	grant_01,
	native_reconfig_writedata_16,
	native_reconfig_writedata_17,
	native_reconfig_writedata_18,
	native_reconfig_writedata_19,
	native_reconfig_writedata_20,
	native_reconfig_writedata_21,
	native_reconfig_writedata_22,
	native_reconfig_writedata_23,
	native_reconfig_writedata_24,
	native_reconfig_writedata_25,
	native_reconfig_writedata_26,
	native_reconfig_writedata_27,
	native_reconfig_writedata_28,
	native_reconfig_writedata_29,
	native_reconfig_writedata_30,
	native_reconfig_writedata_31,
	native_reconfig_write_1,
	native_reconfig_read_1,
	native_reconfig_address_12,
	native_reconfig_address_13,
	native_reconfig_address_14,
	native_reconfig_address_15,
	native_reconfig_address_16,
	native_reconfig_address_17,
	native_reconfig_address_18,
	native_reconfig_address_19,
	native_reconfig_address_20,
	native_reconfig_address_21,
	native_reconfig_address_22,
	native_reconfig_address_23,
	pif_testbus_sel_12,
	pif_testbus_sel_13,
	pif_testbus_sel_14,
	pif_testbus_sel_15,
	reg_plock,
	mutex_grant3,
	mutex_grant4,
	lif_waitrequest1,
	master_read,
	wbasic_read_82,
	lif_waitrequest2,
	basic_reconfig_waitrequest2,
	wbasic_writedata_1_8,
	wbasic_writedata_2_8,
	wbasic_writedata_0_8,
	wbasic_writedata_3_8,
	wbasic_writedata_4_8,
	wbasic_writedata_5_8,
	wbasic_writedata_6_8,
	wbasic_writedata_7_8,
	wbasic_writedata_8_8,
	wbasic_writedata_9_8,
	wbasic_writedata_10_8,
	wbasic_writedata_11_8,
	master_writedata_121,
	master_write_data_12,
	master_writedata_122,
	master_writedata_131,
	master_write_data_13,
	master_writedata_132,
	master_writedata_141,
	master_write_data_14,
	master_writedata_142,
	master_writedata_151,
	master_write_data_15,
	master_writedata_152,
	wbasic_write_83,
	lif_is_active,
	out_narrow_0,
	out_narrow_1,
	out_narrow_2,
	out_narrow_3,
	GND_port,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_16,
	reconfig_from_xcvr_0,
	reconfig_from_xcvr_46,
	reconfig_mgmt_writedata_17,
	reconfig_from_xcvr_1,
	reconfig_from_xcvr_47,
	reconfig_mgmt_writedata_18,
	reconfig_from_xcvr_2,
	reconfig_from_xcvr_48,
	reconfig_mgmt_writedata_19,
	reconfig_from_xcvr_3,
	reconfig_from_xcvr_49,
	reconfig_mgmt_writedata_20,
	reconfig_from_xcvr_4,
	reconfig_from_xcvr_50,
	reconfig_mgmt_writedata_21,
	reconfig_from_xcvr_5,
	reconfig_from_xcvr_51,
	reconfig_mgmt_writedata_22,
	reconfig_from_xcvr_6,
	reconfig_from_xcvr_52,
	reconfig_mgmt_writedata_23,
	reconfig_from_xcvr_7,
	reconfig_from_xcvr_53,
	reconfig_mgmt_writedata_24,
	reconfig_from_xcvr_8,
	reconfig_from_xcvr_54,
	reconfig_mgmt_writedata_25,
	reconfig_from_xcvr_9,
	reconfig_from_xcvr_55,
	reconfig_mgmt_writedata_26,
	reconfig_from_xcvr_10,
	reconfig_from_xcvr_56,
	reconfig_mgmt_writedata_27,
	reconfig_from_xcvr_11,
	reconfig_from_xcvr_57,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_from_xcvr_12,
	reconfig_from_xcvr_58,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_from_xcvr_13,
	reconfig_from_xcvr_59,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_from_xcvr_14,
	reconfig_from_xcvr_60,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15,
	reconfig_from_xcvr_15,
	reconfig_from_xcvr_61,
	reconfig_from_xcvr_24,
	reconfig_from_xcvr_70,
	reconfig_from_xcvr_16,
	reconfig_from_xcvr_62,
	reconfig_from_xcvr_32,
	reconfig_from_xcvr_78,
	reconfig_from_xcvr_25,
	reconfig_from_xcvr_71,
	reconfig_from_xcvr_17,
	reconfig_from_xcvr_63,
	reconfig_from_xcvr_33,
	reconfig_from_xcvr_79,
	reconfig_from_xcvr_26,
	reconfig_from_xcvr_72,
	reconfig_from_xcvr_18,
	reconfig_from_xcvr_64,
	reconfig_from_xcvr_34,
	reconfig_from_xcvr_80,
	reconfig_from_xcvr_27,
	reconfig_from_xcvr_73,
	reconfig_from_xcvr_19,
	reconfig_from_xcvr_65,
	reconfig_from_xcvr_35,
	reconfig_from_xcvr_81)/* synthesis synthesis_greybox=0 */;
output 	basic_reconfig_readdata_12;
output 	basic_reconfig_readdata_13;
output 	basic_reconfig_readdata_14;
output 	basic_reconfig_readdata_15;
output 	basic_reconfig_readdata_16;
output 	basic_reconfig_readdata_17;
output 	basic_reconfig_readdata_18;
output 	basic_reconfig_readdata_19;
output 	basic_reconfig_readdata_20;
output 	basic_reconfig_readdata_21;
output 	basic_reconfig_readdata_22;
output 	basic_reconfig_readdata_23;
output 	basic_reconfig_readdata_24;
output 	basic_reconfig_readdata_25;
output 	basic_reconfig_readdata_26;
output 	basic_reconfig_readdata_27;
output 	basic_reconfig_readdata_28;
output 	basic_reconfig_readdata_29;
output 	basic_reconfig_readdata_30;
output 	basic_reconfig_readdata_31;
input 	master_writedata_16;
input 	master_writedata_17;
input 	master_writedata_18;
input 	master_writedata_19;
input 	master_writedata_20;
input 	master_writedata_21;
input 	master_writedata_22;
input 	master_writedata_23;
input 	master_writedata_24;
input 	master_writedata_25;
input 	master_writedata_26;
input 	master_writedata_27;
input 	master_writedata_28;
input 	master_writedata_12;
input 	master_writedata_29;
input 	master_writedata_13;
input 	master_writedata_30;
input 	master_writedata_14;
input 	master_writedata_31;
input 	master_writedata_15;
output 	basic_reconfig_readdata_0;
output 	basic_reconfig_readdata_1;
output 	basic_reconfig_readdata_2;
output 	basic_reconfig_readdata_3;
output 	basic_reconfig_readdata_4;
output 	basic_reconfig_readdata_5;
input 	Equal2;
output 	basic_reconfig_readdata_6;
output 	basic_reconfig_readdata_7;
output 	basic_reconfig_readdata_8;
output 	basic_reconfig_readdata_9;
output 	basic_reconfig_readdata_10;
output 	basic_reconfig_readdata_11;
input 	mutex_grant;
input 	master_write;
input 	wbasic_write_8;
input 	wbasic_write_81;
input 	wbasic_write_82;
input 	mutex_grant1;
input 	wbasic_address_2_8;
input 	mutex_grant2;
input 	wbasic_address_0_8;
input 	wbasic_address_1_8;
output 	lif_waitrequest;
input 	wbasic_read_8;
input 	wbasic_read_81;
output 	basic_reconfig_waitrequest;
output 	basic_reconfig_waitrequest1;
input 	resync_chains0sync_r_1;
output 	pif_ena_0;
input 	grant_0;
output 	native_reconfig_writedata_0;
output 	native_reconfig_writedata_1;
output 	native_reconfig_writedata_2;
output 	native_reconfig_writedata_3;
output 	native_reconfig_writedata_4;
output 	native_reconfig_writedata_5;
output 	native_reconfig_writedata_6;
output 	native_reconfig_writedata_7;
output 	native_reconfig_writedata_8;
output 	native_reconfig_writedata_9;
output 	native_reconfig_writedata_10;
output 	native_reconfig_writedata_11;
output 	native_reconfig_writedata_12;
output 	native_reconfig_writedata_13;
output 	native_reconfig_writedata_14;
output 	native_reconfig_writedata_15;
output 	native_reconfig_write_0;
output 	native_reconfig_read_0;
output 	native_reconfig_address_0;
output 	native_reconfig_address_1;
output 	native_reconfig_address_2;
output 	native_reconfig_address_3;
output 	native_reconfig_address_4;
output 	native_reconfig_address_5;
output 	native_reconfig_address_6;
output 	native_reconfig_address_7;
output 	native_reconfig_address_8;
output 	native_reconfig_address_9;
output 	native_reconfig_address_10;
output 	native_reconfig_address_11;
output 	pif_testbus_sel_0;
output 	pif_testbus_sel_1;
output 	pif_testbus_sel_2;
output 	pif_testbus_sel_3;
output 	pif_ena_1;
input 	grant_01;
output 	native_reconfig_writedata_16;
output 	native_reconfig_writedata_17;
output 	native_reconfig_writedata_18;
output 	native_reconfig_writedata_19;
output 	native_reconfig_writedata_20;
output 	native_reconfig_writedata_21;
output 	native_reconfig_writedata_22;
output 	native_reconfig_writedata_23;
output 	native_reconfig_writedata_24;
output 	native_reconfig_writedata_25;
output 	native_reconfig_writedata_26;
output 	native_reconfig_writedata_27;
output 	native_reconfig_writedata_28;
output 	native_reconfig_writedata_29;
output 	native_reconfig_writedata_30;
output 	native_reconfig_writedata_31;
output 	native_reconfig_write_1;
output 	native_reconfig_read_1;
output 	native_reconfig_address_12;
output 	native_reconfig_address_13;
output 	native_reconfig_address_14;
output 	native_reconfig_address_15;
output 	native_reconfig_address_16;
output 	native_reconfig_address_17;
output 	native_reconfig_address_18;
output 	native_reconfig_address_19;
output 	native_reconfig_address_20;
output 	native_reconfig_address_21;
output 	native_reconfig_address_22;
output 	native_reconfig_address_23;
output 	pif_testbus_sel_12;
output 	pif_testbus_sel_13;
output 	pif_testbus_sel_14;
output 	pif_testbus_sel_15;
output 	reg_plock;
input 	mutex_grant3;
input 	mutex_grant4;
output 	lif_waitrequest1;
input 	master_read;
input 	wbasic_read_82;
output 	lif_waitrequest2;
output 	basic_reconfig_waitrequest2;
input 	wbasic_writedata_1_8;
input 	wbasic_writedata_2_8;
input 	wbasic_writedata_0_8;
input 	wbasic_writedata_3_8;
input 	wbasic_writedata_4_8;
input 	wbasic_writedata_5_8;
input 	wbasic_writedata_6_8;
input 	wbasic_writedata_7_8;
input 	wbasic_writedata_8_8;
input 	wbasic_writedata_9_8;
input 	wbasic_writedata_10_8;
input 	wbasic_writedata_11_8;
input 	master_writedata_121;
input 	master_write_data_12;
input 	master_writedata_122;
input 	master_writedata_131;
input 	master_write_data_13;
input 	master_writedata_132;
input 	master_writedata_141;
input 	master_write_data_14;
input 	master_writedata_142;
input 	master_writedata_151;
input 	master_write_data_15;
input 	master_writedata_152;
input 	wbasic_write_83;
input 	lif_is_active;
output 	out_narrow_0;
output 	out_narrow_1;
output 	out_narrow_2;
output 	out_narrow_3;
input 	GND_port;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_from_xcvr_0;
input 	reconfig_from_xcvr_46;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_from_xcvr_1;
input 	reconfig_from_xcvr_47;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_from_xcvr_2;
input 	reconfig_from_xcvr_48;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_from_xcvr_3;
input 	reconfig_from_xcvr_49;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_from_xcvr_4;
input 	reconfig_from_xcvr_50;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_from_xcvr_5;
input 	reconfig_from_xcvr_51;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_from_xcvr_6;
input 	reconfig_from_xcvr_52;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_from_xcvr_7;
input 	reconfig_from_xcvr_53;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_from_xcvr_8;
input 	reconfig_from_xcvr_54;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_from_xcvr_9;
input 	reconfig_from_xcvr_55;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_from_xcvr_10;
input 	reconfig_from_xcvr_56;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_from_xcvr_11;
input 	reconfig_from_xcvr_57;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_from_xcvr_12;
input 	reconfig_from_xcvr_58;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_from_xcvr_13;
input 	reconfig_from_xcvr_59;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_from_xcvr_14;
input 	reconfig_from_xcvr_60;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;
input 	reconfig_from_xcvr_15;
input 	reconfig_from_xcvr_61;
input 	reconfig_from_xcvr_24;
input 	reconfig_from_xcvr_70;
input 	reconfig_from_xcvr_16;
input 	reconfig_from_xcvr_62;
input 	reconfig_from_xcvr_32;
input 	reconfig_from_xcvr_78;
input 	reconfig_from_xcvr_25;
input 	reconfig_from_xcvr_71;
input 	reconfig_from_xcvr_17;
input 	reconfig_from_xcvr_63;
input 	reconfig_from_xcvr_33;
input 	reconfig_from_xcvr_79;
input 	reconfig_from_xcvr_26;
input 	reconfig_from_xcvr_72;
input 	reconfig_from_xcvr_18;
input 	reconfig_from_xcvr_64;
input 	reconfig_from_xcvr_34;
input 	reconfig_from_xcvr_80;
input 	reconfig_from_xcvr_27;
input 	reconfig_from_xcvr_73;
input 	reconfig_from_xcvr_19;
input 	reconfig_from_xcvr_65;
input 	reconfig_from_xcvr_35;
input 	reconfig_from_xcvr_81;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lif_csr|reg_rwdata[16]~q ;
wire \lif_csr|reg_rwdata[17]~q ;
wire \lif_csr|reg_rwdata[18]~q ;
wire \lif_csr|reg_rwdata[19]~q ;
wire \lif_csr|reg_rwdata[20]~q ;
wire \lif_csr|reg_rwdata[21]~q ;
wire \lif_csr|reg_rwdata[22]~q ;
wire \lif_csr|reg_rwdata[23]~q ;
wire \lif_csr|reg_rwdata[24]~q ;
wire \lif_csr|reg_rwdata[25]~q ;
wire \lif_csr|reg_rwdata[26]~q ;
wire \lif_csr|reg_rwdata[27]~q ;
wire \lif_csr|reg_rwdata[28]~q ;
wire \lif_csr|reg_rwdata[29]~q ;
wire \lif_csr|reg_rwdata[30]~q ;
wire \lif_csr|reg_rwdata[31]~q ;
wire \lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a0~portadataout ;
wire \lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a1~portadataout ;
wire \lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a2~portadataout ;
wire \lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a3~portadataout ;
wire \lif_csr|reco_read_length_cntr[2]~q ;
wire \lif_csr|reco_read_length_cntr[1]~q ;
wire \lif_csr|reco_read_length_cntr[0]~q ;
wire \lif_csr|reco_addr[11]~q ;
wire \lif_csr|reg_rwdata[0]~q ;
wire \lif_csr|reg_rwdata[1]~q ;
wire \lif_csr|reg_rwdata[2]~q ;
wire \lif_csr|reg_rwdata[3]~q ;
wire \lif_csr|reg_rwdata[4]~q ;
wire \lif_csr|reg_rwdata[5]~q ;
wire \lif_csr|reg_rwdata[6]~q ;
wire \lif_csr|reg_rwdata[7]~q ;
wire \lif_csr|reg_rwdata[8]~q ;
wire \lif_csr|reg_rwdata[9]~q ;
wire \lif_csr|reg_rwdata[10]~q ;
wire \lif_csr|reg_rwdata[11]~q ;
wire \lif_csr|reg_rwdata[12]~q ;
wire \lif_csr|reg_rwdata[13]~q ;
wire \lif_csr|reg_rwdata[14]~q ;
wire \lif_csr|reg_rwdata[15]~q ;
wire \lif_csr|reco_write~q ;
wire \lif_csr|reco_addr[0]~q ;
wire \lif_csr|reco_addr[1]~q ;
wire \lif_csr|reco_addr[2]~q ;
wire \lif_csr|reco_addr[3]~q ;
wire \lif_csr|reco_addr[4]~q ;
wire \lif_csr|reco_addr[5]~q ;
wire \lif_csr|reco_addr[6]~q ;
wire \lif_csr|reco_addr[7]~q ;
wire \lif_csr|reco_addr[8]~q ;
wire \lif_csr|reco_addr[9]~q ;
wire \lif_csr|reco_addr[10]~q ;
wire \lif_csr|testbus_sel[0]~q ;
wire \lif_csr|testbus_sel[1]~q ;
wire \lif_csr|testbus_sel[2]~q ;
wire \lif_csr|testbus_sel[3]~q ;
wire \lif_csr|lif_number[0]~q ;
wire \lif_csr|lif_number[4]~q ;
wire \lif_csr|lif_number[3]~q ;
wire \lif_csr|lif_number[2]~q ;
wire \lif_csr|lif_number[1]~q ;
wire \pif_testbus_groups[1][0]~combout ;
wire \pif_testbus_groups[1][16]~combout ;
wire \pif_testbus_groups[1][1]~combout ;
wire \pif_testbus_groups[1][17]~combout ;
wire \pif_testbus_groups[1][2]~combout ;
wire \pif_testbus_groups[1][18]~combout ;
wire \pif_testbus_groups[1][3]~combout ;
wire \pif_testbus_groups[1][19]~combout ;
wire \pif_ena[0]~0_combout ;
wire \Equal0~0_combout ;
wire \lif_ena[0]~q ;
wire \sel_enabled_and_granted[0]~0_combout ;
wire \upper_16_sel~0_combout ;
wire \upper_16_sel~q ;
wire \pif_enabled_and_granted[0]~combout ;
wire \Equal1~0_combout ;
wire \lif_ena[1]~q ;
wire \sel_enabled_and_granted[1]~1_combout ;
wire \pif_enabled_and_granted[1]~combout ;


RECONFIGURE_IP_csr_mux pif_tbus_mux(
	.ram_block1a0(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a1(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a2(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a2~portadataout ),
	.pif_enabled_and_granted_0(\pif_enabled_and_granted[0]~combout ),
	.pif_enabled_and_granted_1(\pif_enabled_and_granted[1]~combout ),
	.pif_testbus_groups_0_1(\pif_testbus_groups[1][0]~combout ),
	.pif_testbus_groups_16_1(\pif_testbus_groups[1][16]~combout ),
	.out_narrow_0(out_narrow_0),
	.pif_testbus_groups_1_1(\pif_testbus_groups[1][1]~combout ),
	.pif_testbus_groups_17_1(\pif_testbus_groups[1][17]~combout ),
	.out_narrow_1(out_narrow_1),
	.pif_testbus_groups_2_1(\pif_testbus_groups[1][2]~combout ),
	.pif_testbus_groups_18_1(\pif_testbus_groups[1][18]~combout ),
	.out_narrow_2(out_narrow_2),
	.pif_testbus_groups_3_1(\pif_testbus_groups[1][3]~combout ),
	.pif_testbus_groups_19_1(\pif_testbus_groups[1][19]~combout ),
	.out_narrow_3(out_narrow_3),
	.reconfig_from_xcvr_24(reconfig_from_xcvr_24),
	.reconfig_from_xcvr_70(reconfig_from_xcvr_70),
	.reconfig_from_xcvr_25(reconfig_from_xcvr_25),
	.reconfig_from_xcvr_71(reconfig_from_xcvr_71),
	.reconfig_from_xcvr_26(reconfig_from_xcvr_26),
	.reconfig_from_xcvr_72(reconfig_from_xcvr_72),
	.reconfig_from_xcvr_27(reconfig_from_xcvr_27),
	.reconfig_from_xcvr_73(reconfig_from_xcvr_73));

RECONFIGURE_IP_av_xrbasic_lif_csr lif_csr(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.reg_rwdata_16(\lif_csr|reg_rwdata[16]~q ),
	.reg_rwdata_17(\lif_csr|reg_rwdata[17]~q ),
	.reg_rwdata_18(\lif_csr|reg_rwdata[18]~q ),
	.reg_rwdata_19(\lif_csr|reg_rwdata[19]~q ),
	.reg_rwdata_20(\lif_csr|reg_rwdata[20]~q ),
	.reg_rwdata_21(\lif_csr|reg_rwdata[21]~q ),
	.reg_rwdata_22(\lif_csr|reg_rwdata[22]~q ),
	.reg_rwdata_23(\lif_csr|reg_rwdata[23]~q ),
	.reg_rwdata_24(\lif_csr|reg_rwdata[24]~q ),
	.reg_rwdata_25(\lif_csr|reg_rwdata[25]~q ),
	.reg_rwdata_26(\lif_csr|reg_rwdata[26]~q ),
	.reg_rwdata_27(\lif_csr|reg_rwdata[27]~q ),
	.reg_rwdata_28(\lif_csr|reg_rwdata[28]~q ),
	.reg_rwdata_29(\lif_csr|reg_rwdata[29]~q ),
	.reg_rwdata_30(\lif_csr|reg_rwdata[30]~q ),
	.reg_rwdata_31(\lif_csr|reg_rwdata[31]~q ),
	.ram_block1a0(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a1(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a2(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a3(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a3~portadataout ),
	.master_writedata_16(master_writedata_16),
	.master_writedata_17(master_writedata_17),
	.master_writedata_18(master_writedata_18),
	.master_writedata_19(master_writedata_19),
	.master_writedata_20(master_writedata_20),
	.master_writedata_21(master_writedata_21),
	.master_writedata_22(master_writedata_22),
	.master_writedata_23(master_writedata_23),
	.master_writedata_24(master_writedata_24),
	.master_writedata_25(master_writedata_25),
	.master_writedata_26(master_writedata_26),
	.master_writedata_27(master_writedata_27),
	.master_writedata_28(master_writedata_28),
	.master_writedata_12(master_writedata_12),
	.master_writedata_29(master_writedata_29),
	.master_writedata_13(master_writedata_13),
	.master_writedata_30(master_writedata_30),
	.master_writedata_14(master_writedata_14),
	.master_writedata_31(master_writedata_31),
	.master_writedata_15(master_writedata_15),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.Equal2(Equal2),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.mutex_grant(mutex_grant),
	.master_write(master_write),
	.wbasic_write_8(wbasic_write_8),
	.wbasic_write_81(wbasic_write_81),
	.wbasic_write_82(wbasic_write_82),
	.mutex_grant1(mutex_grant1),
	.wbasic_address_2_8(wbasic_address_2_8),
	.mutex_grant2(mutex_grant2),
	.wbasic_address_0_8(wbasic_address_0_8),
	.wbasic_address_1_8(wbasic_address_1_8),
	.lif_waitrequest(lif_waitrequest),
	.wbasic_read_8(wbasic_read_8),
	.wbasic_read_81(wbasic_read_81),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.reco_read_length_cntr_2(\lif_csr|reco_read_length_cntr[2]~q ),
	.reco_read_length_cntr_1(\lif_csr|reco_read_length_cntr[1]~q ),
	.reco_read_length_cntr_0(\lif_csr|reco_read_length_cntr[0]~q ),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.reset(resync_chains0sync_r_1),
	.reco_addr_11(\lif_csr|reco_addr[11]~q ),
	.sel_enabled_and_granted_0(\sel_enabled_and_granted[0]~0_combout ),
	.reg_rwdata_0(\lif_csr|reg_rwdata[0]~q ),
	.reg_rwdata_1(\lif_csr|reg_rwdata[1]~q ),
	.reg_rwdata_2(\lif_csr|reg_rwdata[2]~q ),
	.reg_rwdata_3(\lif_csr|reg_rwdata[3]~q ),
	.reg_rwdata_4(\lif_csr|reg_rwdata[4]~q ),
	.reg_rwdata_5(\lif_csr|reg_rwdata[5]~q ),
	.reg_rwdata_6(\lif_csr|reg_rwdata[6]~q ),
	.reg_rwdata_7(\lif_csr|reg_rwdata[7]~q ),
	.reg_rwdata_8(\lif_csr|reg_rwdata[8]~q ),
	.reg_rwdata_9(\lif_csr|reg_rwdata[9]~q ),
	.reg_rwdata_10(\lif_csr|reg_rwdata[10]~q ),
	.reg_rwdata_11(\lif_csr|reg_rwdata[11]~q ),
	.reg_rwdata_12(\lif_csr|reg_rwdata[12]~q ),
	.reg_rwdata_13(\lif_csr|reg_rwdata[13]~q ),
	.reg_rwdata_14(\lif_csr|reg_rwdata[14]~q ),
	.reg_rwdata_15(\lif_csr|reg_rwdata[15]~q ),
	.reco_write1(\lif_csr|reco_write~q ),
	.reco_addr_0(\lif_csr|reco_addr[0]~q ),
	.reco_addr_1(\lif_csr|reco_addr[1]~q ),
	.reco_addr_2(\lif_csr|reco_addr[2]~q ),
	.reco_addr_3(\lif_csr|reco_addr[3]~q ),
	.reco_addr_4(\lif_csr|reco_addr[4]~q ),
	.reco_addr_5(\lif_csr|reco_addr[5]~q ),
	.reco_addr_6(\lif_csr|reco_addr[6]~q ),
	.reco_addr_7(\lif_csr|reco_addr[7]~q ),
	.reco_addr_8(\lif_csr|reco_addr[8]~q ),
	.reco_addr_9(\lif_csr|reco_addr[9]~q ),
	.reco_addr_10(\lif_csr|reco_addr[10]~q ),
	.pif_enabled_and_granted_0(\pif_enabled_and_granted[0]~combout ),
	.testbus_sel_0(\lif_csr|testbus_sel[0]~q ),
	.testbus_sel_1(\lif_csr|testbus_sel[1]~q ),
	.testbus_sel_2(\lif_csr|testbus_sel[2]~q ),
	.testbus_sel_3(\lif_csr|testbus_sel[3]~q ),
	.sel_enabled_and_granted_1(\sel_enabled_and_granted[1]~1_combout ),
	.pif_enabled_and_granted_1(\pif_enabled_and_granted[1]~combout ),
	.reg_plock1(reg_plock),
	.mutex_grant3(mutex_grant3),
	.mutex_grant4(mutex_grant4),
	.lif_waitrequest1(lif_waitrequest1),
	.master_read(master_read),
	.wbasic_read_82(wbasic_read_82),
	.lif_waitrequest2(lif_waitrequest2),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.wbasic_writedata_1_8(wbasic_writedata_1_8),
	.wbasic_writedata_2_8(wbasic_writedata_2_8),
	.wbasic_writedata_0_8(wbasic_writedata_0_8),
	.wbasic_writedata_3_8(wbasic_writedata_3_8),
	.lif_number_0(\lif_csr|lif_number[0]~q ),
	.lif_number_4(\lif_csr|lif_number[4]~q ),
	.lif_number_3(\lif_csr|lif_number[3]~q ),
	.lif_number_2(\lif_csr|lif_number[2]~q ),
	.lif_number_1(\lif_csr|lif_number[1]~q ),
	.wbasic_writedata_4_8(wbasic_writedata_4_8),
	.wbasic_writedata_5_8(wbasic_writedata_5_8),
	.wbasic_writedata_6_8(wbasic_writedata_6_8),
	.wbasic_writedata_7_8(wbasic_writedata_7_8),
	.wbasic_writedata_8_8(wbasic_writedata_8_8),
	.wbasic_writedata_9_8(wbasic_writedata_9_8),
	.wbasic_writedata_10_8(wbasic_writedata_10_8),
	.wbasic_writedata_11_8(wbasic_writedata_11_8),
	.master_writedata_121(master_writedata_121),
	.master_write_data_12(master_write_data_12),
	.master_writedata_122(master_writedata_122),
	.master_writedata_131(master_writedata_131),
	.master_write_data_13(master_write_data_13),
	.master_writedata_132(master_writedata_132),
	.master_writedata_141(master_writedata_141),
	.master_write_data_14(master_write_data_14),
	.master_writedata_142(master_writedata_142),
	.master_writedata_151(master_writedata_151),
	.master_write_data_15(master_write_data_15),
	.master_writedata_152(master_writedata_152),
	.wbasic_write_83(wbasic_write_83),
	.lif_is_active(lif_is_active),
	.GND_port(GND_port),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_from_xcvr_0(reconfig_from_xcvr_0),
	.reconfig_from_xcvr_46(reconfig_from_xcvr_46),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_from_xcvr_1(reconfig_from_xcvr_1),
	.reconfig_from_xcvr_47(reconfig_from_xcvr_47),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_from_xcvr_2(reconfig_from_xcvr_2),
	.reconfig_from_xcvr_48(reconfig_from_xcvr_48),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_from_xcvr_3(reconfig_from_xcvr_3),
	.reconfig_from_xcvr_49(reconfig_from_xcvr_49),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_from_xcvr_4(reconfig_from_xcvr_4),
	.reconfig_from_xcvr_50(reconfig_from_xcvr_50),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_from_xcvr_5(reconfig_from_xcvr_5),
	.reconfig_from_xcvr_51(reconfig_from_xcvr_51),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_from_xcvr_6(reconfig_from_xcvr_6),
	.reconfig_from_xcvr_52(reconfig_from_xcvr_52),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_from_xcvr_7(reconfig_from_xcvr_7),
	.reconfig_from_xcvr_53(reconfig_from_xcvr_53),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_from_xcvr_8(reconfig_from_xcvr_8),
	.reconfig_from_xcvr_54(reconfig_from_xcvr_54),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_from_xcvr_9(reconfig_from_xcvr_9),
	.reconfig_from_xcvr_55(reconfig_from_xcvr_55),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_from_xcvr_10(reconfig_from_xcvr_10),
	.reconfig_from_xcvr_56(reconfig_from_xcvr_56),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_from_xcvr_11(reconfig_from_xcvr_11),
	.reconfig_from_xcvr_57(reconfig_from_xcvr_57),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_from_xcvr_12(reconfig_from_xcvr_12),
	.reconfig_from_xcvr_58(reconfig_from_xcvr_58),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_from_xcvr_13(reconfig_from_xcvr_13),
	.reconfig_from_xcvr_59(reconfig_from_xcvr_59),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_from_xcvr_14(reconfig_from_xcvr_14),
	.reconfig_from_xcvr_60(reconfig_from_xcvr_60),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15),
	.reconfig_from_xcvr_15(reconfig_from_xcvr_15),
	.reconfig_from_xcvr_61(reconfig_from_xcvr_61));

cyclonev_lcell_comb \pif_testbus_groups[1][0] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_16),
	.dataf(!reconfig_from_xcvr_62),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][0] .extended_lut = "off";
defparam \pif_testbus_groups[1][0] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][0] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_groups[1][16] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_32),
	.dataf(!reconfig_from_xcvr_78),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][16] .extended_lut = "off";
defparam \pif_testbus_groups[1][16] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][16] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_groups[1][1] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_17),
	.dataf(!reconfig_from_xcvr_63),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][1] .extended_lut = "off";
defparam \pif_testbus_groups[1][1] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][1] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_groups[1][17] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_33),
	.dataf(!reconfig_from_xcvr_79),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][17] .extended_lut = "off";
defparam \pif_testbus_groups[1][17] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][17] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_groups[1][2] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_18),
	.dataf(!reconfig_from_xcvr_64),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][2] .extended_lut = "off";
defparam \pif_testbus_groups[1][2] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][2] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_groups[1][18] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_34),
	.dataf(!reconfig_from_xcvr_80),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][18] .extended_lut = "off";
defparam \pif_testbus_groups[1][18] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][18] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_groups[1][3] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_19),
	.dataf(!reconfig_from_xcvr_65),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][3] .extended_lut = "off";
defparam \pif_testbus_groups[1][3] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][3] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_groups[1][19] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(!reconfig_from_xcvr_35),
	.dataf(!reconfig_from_xcvr_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_testbus_groups[1][19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_groups[1][19] .extended_lut = "off";
defparam \pif_testbus_groups[1][19] .lut_mask = 64'h00001111000F111F;
defparam \pif_testbus_groups[1][19] .shared_arith = "off";

dffeas \pif_ena[0] (
	.clk(mgmt_clk_clk),
	.d(\pif_ena[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pif_ena_0),
	.prn(vcc));
defparam \pif_ena[0] .is_wysiwyg = "true";
defparam \pif_ena[0] .power_up = "low";

cyclonev_lcell_comb \native_reconfig_writedata[0]~0 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[16]~q ),
	.datad(!\lif_csr|reg_rwdata[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[0]~0 .extended_lut = "off";
defparam \native_reconfig_writedata[0]~0 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[1]~1 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[17]~q ),
	.datad(!\lif_csr|reg_rwdata[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[1]~1 .extended_lut = "off";
defparam \native_reconfig_writedata[1]~1 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[2]~2 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[18]~q ),
	.datad(!\lif_csr|reg_rwdata[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[2]~2 .extended_lut = "off";
defparam \native_reconfig_writedata[2]~2 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[3]~3 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[19]~q ),
	.datad(!\lif_csr|reg_rwdata[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[3]~3 .extended_lut = "off";
defparam \native_reconfig_writedata[3]~3 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[4]~4 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[20]~q ),
	.datad(!\lif_csr|reg_rwdata[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[4]~4 .extended_lut = "off";
defparam \native_reconfig_writedata[4]~4 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[5]~5 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[21]~q ),
	.datad(!\lif_csr|reg_rwdata[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[5]~5 .extended_lut = "off";
defparam \native_reconfig_writedata[5]~5 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[6]~6 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[22]~q ),
	.datad(!\lif_csr|reg_rwdata[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[6]~6 .extended_lut = "off";
defparam \native_reconfig_writedata[6]~6 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[7]~7 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[23]~q ),
	.datad(!\lif_csr|reg_rwdata[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[7]~7 .extended_lut = "off";
defparam \native_reconfig_writedata[7]~7 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[8]~8 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[24]~q ),
	.datad(!\lif_csr|reg_rwdata[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[8]~8 .extended_lut = "off";
defparam \native_reconfig_writedata[8]~8 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[9]~9 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[25]~q ),
	.datad(!\lif_csr|reg_rwdata[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[9]~9 .extended_lut = "off";
defparam \native_reconfig_writedata[9]~9 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[9]~9 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[10]~10 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[26]~q ),
	.datad(!\lif_csr|reg_rwdata[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[10]~10 .extended_lut = "off";
defparam \native_reconfig_writedata[10]~10 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[10]~10 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[11]~11 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[27]~q ),
	.datad(!\lif_csr|reg_rwdata[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[11]~11 .extended_lut = "off";
defparam \native_reconfig_writedata[11]~11 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[11]~11 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[12]~12 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[28]~q ),
	.datad(!\lif_csr|reg_rwdata[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[12]~12 .extended_lut = "off";
defparam \native_reconfig_writedata[12]~12 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[12]~12 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[13]~13 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[29]~q ),
	.datad(!\lif_csr|reg_rwdata[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[13]~13 .extended_lut = "off";
defparam \native_reconfig_writedata[13]~13 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[13]~13 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[14]~14 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[30]~q ),
	.datad(!\lif_csr|reg_rwdata[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[14]~14 .extended_lut = "off";
defparam \native_reconfig_writedata[14]~14 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[14]~14 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[15]~15 (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\upper_16_sel~q ),
	.datac(!\lif_csr|reg_rwdata[31]~q ),
	.datad(!\lif_csr|reg_rwdata[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[15]~15 .extended_lut = "off";
defparam \native_reconfig_writedata[15]~15 .lut_mask = 64'h0145014501450145;
defparam \native_reconfig_writedata[15]~15 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_write[0] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_write~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_write_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_write[0] .extended_lut = "off";
defparam \native_reconfig_write[0] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_write[0] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_read[0]~0 (
	.dataa(!\lif_csr|reco_read_length_cntr[2]~q ),
	.datab(!\lif_csr|reco_read_length_cntr[1]~q ),
	.datac(!\lif_csr|reco_read_length_cntr[0]~q ),
	.datad(!\sel_enabled_and_granted[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_read_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_read[0]~0 .extended_lut = "off";
defparam \native_reconfig_read[0]~0 .lut_mask = 64'h0057005700570057;
defparam \native_reconfig_read[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[0] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[0] .extended_lut = "off";
defparam \native_reconfig_address[0] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[0] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[1] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[1] .extended_lut = "off";
defparam \native_reconfig_address[1] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[1] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[2] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[2] .extended_lut = "off";
defparam \native_reconfig_address[2] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[2] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[3] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[3] .extended_lut = "off";
defparam \native_reconfig_address[3] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[3] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[4] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[4] .extended_lut = "off";
defparam \native_reconfig_address[4] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[4] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[5] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[5] .extended_lut = "off";
defparam \native_reconfig_address[5] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[5] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[6] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[6] .extended_lut = "off";
defparam \native_reconfig_address[6] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[6] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[7] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[7] .extended_lut = "off";
defparam \native_reconfig_address[7] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[7] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[8] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[8] .extended_lut = "off";
defparam \native_reconfig_address[8] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[8] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[9] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[9] .extended_lut = "off";
defparam \native_reconfig_address[9] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[9] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[10] (
	.dataa(!\sel_enabled_and_granted[0]~0_combout ),
	.datab(!\lif_csr|reco_addr[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[10] .extended_lut = "off";
defparam \native_reconfig_address[10] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[10] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[11]~0 (
	.dataa(!\lif_ena[0]~q ),
	.datab(!\lif_csr|reco_addr[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[11]~0 .extended_lut = "off";
defparam \native_reconfig_address[11]~0 .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[11]~0 .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[0] (
	.dataa(!\pif_enabled_and_granted[0]~combout ),
	.datab(!\lif_csr|testbus_sel[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[0] .extended_lut = "off";
defparam \pif_testbus_sel[0] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[0] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[1] (
	.dataa(!\pif_enabled_and_granted[0]~combout ),
	.datab(!\lif_csr|testbus_sel[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[1] .extended_lut = "off";
defparam \pif_testbus_sel[1] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[1] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[2] (
	.dataa(!\pif_enabled_and_granted[0]~combout ),
	.datab(!\lif_csr|testbus_sel[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[2] .extended_lut = "off";
defparam \pif_testbus_sel[2] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[2] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[3] (
	.dataa(!\pif_enabled_and_granted[0]~combout ),
	.datab(!\lif_csr|testbus_sel[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[3] .extended_lut = "off";
defparam \pif_testbus_sel[3] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[3] .shared_arith = "off";

dffeas \pif_ena[1] (
	.clk(mgmt_clk_clk),
	.d(\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a3~portadataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pif_ena_1),
	.prn(vcc));
defparam \pif_ena[1] .is_wysiwyg = "true";
defparam \pif_ena[1] .power_up = "low";

cyclonev_lcell_comb \native_reconfig_writedata[16]~16 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[16]~q ),
	.datac(!\lif_csr|reg_rwdata[0]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[16]~16 .extended_lut = "off";
defparam \native_reconfig_writedata[16]~16 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[16]~16 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[17]~17 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[17]~q ),
	.datac(!\lif_csr|reg_rwdata[1]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[17]~17 .extended_lut = "off";
defparam \native_reconfig_writedata[17]~17 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[17]~17 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[18]~18 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[18]~q ),
	.datac(!\lif_csr|reg_rwdata[2]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[18]~18 .extended_lut = "off";
defparam \native_reconfig_writedata[18]~18 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[18]~18 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[19]~19 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[19]~q ),
	.datac(!\lif_csr|reg_rwdata[3]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[19]~19 .extended_lut = "off";
defparam \native_reconfig_writedata[19]~19 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[19]~19 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[20]~20 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[20]~q ),
	.datac(!\lif_csr|reg_rwdata[4]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[20]~20 .extended_lut = "off";
defparam \native_reconfig_writedata[20]~20 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[20]~20 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[21]~21 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[21]~q ),
	.datac(!\lif_csr|reg_rwdata[5]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[21]~21 .extended_lut = "off";
defparam \native_reconfig_writedata[21]~21 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[21]~21 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[22]~22 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[22]~q ),
	.datac(!\lif_csr|reg_rwdata[6]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[22]~22 .extended_lut = "off";
defparam \native_reconfig_writedata[22]~22 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[22]~22 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[23]~23 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[23]~q ),
	.datac(!\lif_csr|reg_rwdata[7]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[23]~23 .extended_lut = "off";
defparam \native_reconfig_writedata[23]~23 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[23]~23 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[24]~24 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[24]~q ),
	.datac(!\lif_csr|reg_rwdata[8]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[24]~24 .extended_lut = "off";
defparam \native_reconfig_writedata[24]~24 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[24]~24 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[25]~25 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[25]~q ),
	.datac(!\lif_csr|reg_rwdata[9]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[25]~25 .extended_lut = "off";
defparam \native_reconfig_writedata[25]~25 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[25]~25 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[26]~26 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[26]~q ),
	.datac(!\lif_csr|reg_rwdata[10]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[26]~26 .extended_lut = "off";
defparam \native_reconfig_writedata[26]~26 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[26]~26 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[27]~27 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[27]~q ),
	.datac(!\lif_csr|reg_rwdata[11]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[27]~27 .extended_lut = "off";
defparam \native_reconfig_writedata[27]~27 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[27]~27 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[28]~28 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[28]~q ),
	.datac(!\lif_csr|reg_rwdata[12]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[28]~28 .extended_lut = "off";
defparam \native_reconfig_writedata[28]~28 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[28]~28 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[29]~29 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[29]~q ),
	.datac(!\lif_csr|reg_rwdata[13]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[29]~29 .extended_lut = "off";
defparam \native_reconfig_writedata[29]~29 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[29]~29 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[30]~30 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[30]~q ),
	.datac(!\lif_csr|reg_rwdata[14]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[30]~30 .extended_lut = "off";
defparam \native_reconfig_writedata[30]~30 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[30]~30 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_writedata[31]~31 (
	.dataa(!\upper_16_sel~q ),
	.datab(!\lif_csr|reg_rwdata[31]~q ),
	.datac(!\lif_csr|reg_rwdata[15]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_writedata_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_writedata[31]~31 .extended_lut = "off";
defparam \native_reconfig_writedata[31]~31 .lut_mask = 64'h001B001B001B001B;
defparam \native_reconfig_writedata[31]~31 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_write[1] (
	.dataa(!\lif_csr|reco_write~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_write_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_write[1] .extended_lut = "off";
defparam \native_reconfig_write[1] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_write[1] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_read[1]~1 (
	.dataa(!\lif_csr|reco_read_length_cntr[2]~q ),
	.datab(!\lif_csr|reco_read_length_cntr[1]~q ),
	.datac(!\lif_csr|reco_read_length_cntr[0]~q ),
	.datad(!\sel_enabled_and_granted[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_read_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_read[1]~1 .extended_lut = "off";
defparam \native_reconfig_read[1]~1 .lut_mask = 64'h0057005700570057;
defparam \native_reconfig_read[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[12] (
	.dataa(!\lif_csr|reco_addr[0]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[12] .extended_lut = "off";
defparam \native_reconfig_address[12] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[12] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[13] (
	.dataa(!\lif_csr|reco_addr[1]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[13] .extended_lut = "off";
defparam \native_reconfig_address[13] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[13] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[14] (
	.dataa(!\lif_csr|reco_addr[2]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[14] .extended_lut = "off";
defparam \native_reconfig_address[14] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[14] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[15] (
	.dataa(!\lif_csr|reco_addr[3]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[15] .extended_lut = "off";
defparam \native_reconfig_address[15] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[15] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[16] (
	.dataa(!\lif_csr|reco_addr[4]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[16] .extended_lut = "off";
defparam \native_reconfig_address[16] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[16] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[17] (
	.dataa(!\lif_csr|reco_addr[5]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[17] .extended_lut = "off";
defparam \native_reconfig_address[17] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[17] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[18] (
	.dataa(!\lif_csr|reco_addr[6]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[18] .extended_lut = "off";
defparam \native_reconfig_address[18] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[18] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[19] (
	.dataa(!\lif_csr|reco_addr[7]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[19] .extended_lut = "off";
defparam \native_reconfig_address[19] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[19] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[20] (
	.dataa(!\lif_csr|reco_addr[8]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[20] .extended_lut = "off";
defparam \native_reconfig_address[20] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[20] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[21] (
	.dataa(!\lif_csr|reco_addr[9]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[21] .extended_lut = "off";
defparam \native_reconfig_address[21] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[21] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[22] (
	.dataa(!\lif_csr|reco_addr[10]~q ),
	.datab(!\sel_enabled_and_granted[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[22] .extended_lut = "off";
defparam \native_reconfig_address[22] .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[22] .shared_arith = "off";

cyclonev_lcell_comb \native_reconfig_address[23]~1 (
	.dataa(!\lif_csr|reco_addr[11]~q ),
	.datab(!\lif_ena[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(native_reconfig_address_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \native_reconfig_address[23]~1 .extended_lut = "off";
defparam \native_reconfig_address[23]~1 .lut_mask = 64'h1111111111111111;
defparam \native_reconfig_address[23]~1 .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[12] (
	.dataa(!\lif_csr|testbus_sel[0]~q ),
	.datab(!\pif_enabled_and_granted[1]~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[12] .extended_lut = "off";
defparam \pif_testbus_sel[12] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[12] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[13] (
	.dataa(!\lif_csr|testbus_sel[1]~q ),
	.datab(!\pif_enabled_and_granted[1]~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[13] .extended_lut = "off";
defparam \pif_testbus_sel[13] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[13] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[14] (
	.dataa(!\lif_csr|testbus_sel[2]~q ),
	.datab(!\pif_enabled_and_granted[1]~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[14] .extended_lut = "off";
defparam \pif_testbus_sel[14] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[14] .shared_arith = "off";

cyclonev_lcell_comb \pif_testbus_sel[15] (
	.dataa(!\lif_csr|testbus_sel[3]~q ),
	.datab(!\pif_enabled_and_granted[1]~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(pif_testbus_sel_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_testbus_sel[15] .extended_lut = "off";
defparam \pif_testbus_sel[15] .lut_mask = 64'h1111111111111111;
defparam \pif_testbus_sel[15] .shared_arith = "off";

cyclonev_lcell_comb \pif_ena[0]~0 (
	.dataa(!\lif_csr|l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a3~portadataout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_ena[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_ena[0]~0 .extended_lut = "off";
defparam \pif_ena[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pif_ena[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\lif_csr|lif_number[0]~q ),
	.datab(!\lif_csr|lif_number[4]~q ),
	.datac(!\lif_csr|lif_number[3]~q ),
	.datad(!\lif_csr|lif_number[2]~q ),
	.datae(!\lif_csr|lif_number[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h8000000080000000;
defparam \Equal0~0 .shared_arith = "off";

dffeas \lif_ena[0] (
	.clk(mgmt_clk_clk),
	.d(\Equal0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lif_ena[0]~q ),
	.prn(vcc));
defparam \lif_ena[0] .is_wysiwyg = "true";
defparam \lif_ena[0] .power_up = "low";

cyclonev_lcell_comb \sel_enabled_and_granted[0]~0 (
	.dataa(!\lif_ena[0]~q ),
	.datab(!\lif_csr|reco_addr[11]~q ),
	.datac(!pif_ena_0),
	.datad(!grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sel_enabled_and_granted[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sel_enabled_and_granted[0]~0 .extended_lut = "off";
defparam \sel_enabled_and_granted[0]~0 .lut_mask = 64'h111D111D111D111D;
defparam \sel_enabled_and_granted[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \upper_16_sel~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\upper_16_sel~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \upper_16_sel~0 .extended_lut = "off";
defparam \upper_16_sel~0 .lut_mask = 64'h0000000000000000;
defparam \upper_16_sel~0 .shared_arith = "off";

dffeas upper_16_sel(
	.clk(mgmt_clk_clk),
	.d(\upper_16_sel~0_combout ),
	.asdata(vcc),
	.clrn(resync_chains0sync_r_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\upper_16_sel~q ),
	.prn(vcc));
defparam upper_16_sel.is_wysiwyg = "true";
defparam upper_16_sel.power_up = "low";

cyclonev_lcell_comb \pif_enabled_and_granted[0] (
	.dataa(!pif_ena_0),
	.datab(!grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_enabled_and_granted[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_enabled_and_granted[0] .extended_lut = "off";
defparam \pif_enabled_and_granted[0] .lut_mask = 64'h1111111111111111;
defparam \pif_enabled_and_granted[0] .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!\lif_csr|lif_number[0]~q ),
	.datab(!\lif_csr|lif_number[4]~q ),
	.datac(!\lif_csr|lif_number[3]~q ),
	.datad(!\lif_csr|lif_number[2]~q ),
	.datae(!\lif_csr|lif_number[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h4000000040000000;
defparam \Equal1~0 .shared_arith = "off";

dffeas \lif_ena[1] (
	.clk(mgmt_clk_clk),
	.d(\Equal1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lif_ena[1]~q ),
	.prn(vcc));
defparam \lif_ena[1] .is_wysiwyg = "true";
defparam \lif_ena[1] .power_up = "low";

cyclonev_lcell_comb \sel_enabled_and_granted[1]~1 (
	.dataa(!\lif_csr|reco_addr[11]~q ),
	.datab(!\lif_ena[1]~q ),
	.datac(!pif_ena_1),
	.datad(!grant_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sel_enabled_and_granted[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sel_enabled_and_granted[1]~1 .extended_lut = "off";
defparam \sel_enabled_and_granted[1]~1 .lut_mask = 64'h111B111B111B111B;
defparam \sel_enabled_and_granted[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \pif_enabled_and_granted[1] (
	.dataa(!pif_ena_1),
	.datab(!grant_01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pif_enabled_and_granted[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pif_enabled_and_granted[1] .extended_lut = "off";
defparam \pif_enabled_and_granted[1] .lut_mask = 64'h1111111111111111;
defparam \pif_enabled_and_granted[1] .shared_arith = "off";

endmodule

module RECONFIGURE_IP_av_xrbasic_lif_csr (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	reg_rwdata_16,
	reg_rwdata_17,
	reg_rwdata_18,
	reg_rwdata_19,
	reg_rwdata_20,
	reg_rwdata_21,
	reg_rwdata_22,
	reg_rwdata_23,
	reg_rwdata_24,
	reg_rwdata_25,
	reg_rwdata_26,
	reg_rwdata_27,
	reg_rwdata_28,
	reg_rwdata_29,
	reg_rwdata_30,
	reg_rwdata_31,
	ram_block1a0,
	ram_block1a1,
	ram_block1a2,
	ram_block1a3,
	master_writedata_16,
	master_writedata_17,
	master_writedata_18,
	master_writedata_19,
	master_writedata_20,
	master_writedata_21,
	master_writedata_22,
	master_writedata_23,
	master_writedata_24,
	master_writedata_25,
	master_writedata_26,
	master_writedata_27,
	master_writedata_28,
	master_writedata_12,
	master_writedata_29,
	master_writedata_13,
	master_writedata_30,
	master_writedata_14,
	master_writedata_31,
	master_writedata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	Equal2,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	mutex_grant,
	master_write,
	wbasic_write_8,
	wbasic_write_81,
	wbasic_write_82,
	mutex_grant1,
	wbasic_address_2_8,
	mutex_grant2,
	wbasic_address_0_8,
	wbasic_address_1_8,
	lif_waitrequest,
	wbasic_read_8,
	wbasic_read_81,
	basic_reconfig_waitrequest,
	reco_read_length_cntr_2,
	reco_read_length_cntr_1,
	reco_read_length_cntr_0,
	basic_reconfig_waitrequest1,
	reset,
	reco_addr_11,
	sel_enabled_and_granted_0,
	reg_rwdata_0,
	reg_rwdata_1,
	reg_rwdata_2,
	reg_rwdata_3,
	reg_rwdata_4,
	reg_rwdata_5,
	reg_rwdata_6,
	reg_rwdata_7,
	reg_rwdata_8,
	reg_rwdata_9,
	reg_rwdata_10,
	reg_rwdata_11,
	reg_rwdata_12,
	reg_rwdata_13,
	reg_rwdata_14,
	reg_rwdata_15,
	reco_write1,
	reco_addr_0,
	reco_addr_1,
	reco_addr_2,
	reco_addr_3,
	reco_addr_4,
	reco_addr_5,
	reco_addr_6,
	reco_addr_7,
	reco_addr_8,
	reco_addr_9,
	reco_addr_10,
	pif_enabled_and_granted_0,
	testbus_sel_0,
	testbus_sel_1,
	testbus_sel_2,
	testbus_sel_3,
	sel_enabled_and_granted_1,
	pif_enabled_and_granted_1,
	reg_plock1,
	mutex_grant3,
	mutex_grant4,
	lif_waitrequest1,
	master_read,
	wbasic_read_82,
	lif_waitrequest2,
	basic_reconfig_waitrequest2,
	wbasic_writedata_1_8,
	wbasic_writedata_2_8,
	wbasic_writedata_0_8,
	wbasic_writedata_3_8,
	lif_number_0,
	lif_number_4,
	lif_number_3,
	lif_number_2,
	lif_number_1,
	wbasic_writedata_4_8,
	wbasic_writedata_5_8,
	wbasic_writedata_6_8,
	wbasic_writedata_7_8,
	wbasic_writedata_8_8,
	wbasic_writedata_9_8,
	wbasic_writedata_10_8,
	wbasic_writedata_11_8,
	master_writedata_121,
	master_write_data_12,
	master_writedata_122,
	master_writedata_131,
	master_write_data_13,
	master_writedata_132,
	master_writedata_141,
	master_write_data_14,
	master_writedata_142,
	master_writedata_151,
	master_write_data_15,
	master_writedata_152,
	wbasic_write_83,
	lif_is_active,
	GND_port,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_16,
	reconfig_from_xcvr_0,
	reconfig_from_xcvr_46,
	reconfig_mgmt_writedata_17,
	reconfig_from_xcvr_1,
	reconfig_from_xcvr_47,
	reconfig_mgmt_writedata_18,
	reconfig_from_xcvr_2,
	reconfig_from_xcvr_48,
	reconfig_mgmt_writedata_19,
	reconfig_from_xcvr_3,
	reconfig_from_xcvr_49,
	reconfig_mgmt_writedata_20,
	reconfig_from_xcvr_4,
	reconfig_from_xcvr_50,
	reconfig_mgmt_writedata_21,
	reconfig_from_xcvr_5,
	reconfig_from_xcvr_51,
	reconfig_mgmt_writedata_22,
	reconfig_from_xcvr_6,
	reconfig_from_xcvr_52,
	reconfig_mgmt_writedata_23,
	reconfig_from_xcvr_7,
	reconfig_from_xcvr_53,
	reconfig_mgmt_writedata_24,
	reconfig_from_xcvr_8,
	reconfig_from_xcvr_54,
	reconfig_mgmt_writedata_25,
	reconfig_from_xcvr_9,
	reconfig_from_xcvr_55,
	reconfig_mgmt_writedata_26,
	reconfig_from_xcvr_10,
	reconfig_from_xcvr_56,
	reconfig_mgmt_writedata_27,
	reconfig_from_xcvr_11,
	reconfig_from_xcvr_57,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_from_xcvr_12,
	reconfig_from_xcvr_58,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_from_xcvr_13,
	reconfig_from_xcvr_59,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_from_xcvr_14,
	reconfig_from_xcvr_60,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15,
	reconfig_from_xcvr_15,
	reconfig_from_xcvr_61)/* synthesis synthesis_greybox=0 */;
output 	basic_reconfig_readdata_12;
output 	basic_reconfig_readdata_13;
output 	basic_reconfig_readdata_14;
output 	basic_reconfig_readdata_15;
output 	basic_reconfig_readdata_16;
output 	basic_reconfig_readdata_17;
output 	basic_reconfig_readdata_18;
output 	basic_reconfig_readdata_19;
output 	basic_reconfig_readdata_20;
output 	basic_reconfig_readdata_21;
output 	basic_reconfig_readdata_22;
output 	basic_reconfig_readdata_23;
output 	basic_reconfig_readdata_24;
output 	basic_reconfig_readdata_25;
output 	basic_reconfig_readdata_26;
output 	basic_reconfig_readdata_27;
output 	basic_reconfig_readdata_28;
output 	basic_reconfig_readdata_29;
output 	basic_reconfig_readdata_30;
output 	basic_reconfig_readdata_31;
output 	reg_rwdata_16;
output 	reg_rwdata_17;
output 	reg_rwdata_18;
output 	reg_rwdata_19;
output 	reg_rwdata_20;
output 	reg_rwdata_21;
output 	reg_rwdata_22;
output 	reg_rwdata_23;
output 	reg_rwdata_24;
output 	reg_rwdata_25;
output 	reg_rwdata_26;
output 	reg_rwdata_27;
output 	reg_rwdata_28;
output 	reg_rwdata_29;
output 	reg_rwdata_30;
output 	reg_rwdata_31;
output 	ram_block1a0;
output 	ram_block1a1;
output 	ram_block1a2;
output 	ram_block1a3;
input 	master_writedata_16;
input 	master_writedata_17;
input 	master_writedata_18;
input 	master_writedata_19;
input 	master_writedata_20;
input 	master_writedata_21;
input 	master_writedata_22;
input 	master_writedata_23;
input 	master_writedata_24;
input 	master_writedata_25;
input 	master_writedata_26;
input 	master_writedata_27;
input 	master_writedata_28;
input 	master_writedata_12;
input 	master_writedata_29;
input 	master_writedata_13;
input 	master_writedata_30;
input 	master_writedata_14;
input 	master_writedata_31;
input 	master_writedata_15;
output 	basic_reconfig_readdata_0;
output 	basic_reconfig_readdata_1;
output 	basic_reconfig_readdata_2;
output 	basic_reconfig_readdata_3;
output 	basic_reconfig_readdata_4;
output 	basic_reconfig_readdata_5;
input 	Equal2;
output 	basic_reconfig_readdata_6;
output 	basic_reconfig_readdata_7;
output 	basic_reconfig_readdata_8;
output 	basic_reconfig_readdata_9;
output 	basic_reconfig_readdata_10;
output 	basic_reconfig_readdata_11;
input 	mutex_grant;
input 	master_write;
input 	wbasic_write_8;
input 	wbasic_write_81;
input 	wbasic_write_82;
input 	mutex_grant1;
input 	wbasic_address_2_8;
input 	mutex_grant2;
input 	wbasic_address_0_8;
input 	wbasic_address_1_8;
output 	lif_waitrequest;
input 	wbasic_read_8;
input 	wbasic_read_81;
output 	basic_reconfig_waitrequest;
output 	reco_read_length_cntr_2;
output 	reco_read_length_cntr_1;
output 	reco_read_length_cntr_0;
output 	basic_reconfig_waitrequest1;
input 	reset;
output 	reco_addr_11;
input 	sel_enabled_and_granted_0;
output 	reg_rwdata_0;
output 	reg_rwdata_1;
output 	reg_rwdata_2;
output 	reg_rwdata_3;
output 	reg_rwdata_4;
output 	reg_rwdata_5;
output 	reg_rwdata_6;
output 	reg_rwdata_7;
output 	reg_rwdata_8;
output 	reg_rwdata_9;
output 	reg_rwdata_10;
output 	reg_rwdata_11;
output 	reg_rwdata_12;
output 	reg_rwdata_13;
output 	reg_rwdata_14;
output 	reg_rwdata_15;
output 	reco_write1;
output 	reco_addr_0;
output 	reco_addr_1;
output 	reco_addr_2;
output 	reco_addr_3;
output 	reco_addr_4;
output 	reco_addr_5;
output 	reco_addr_6;
output 	reco_addr_7;
output 	reco_addr_8;
output 	reco_addr_9;
output 	reco_addr_10;
input 	pif_enabled_and_granted_0;
output 	testbus_sel_0;
output 	testbus_sel_1;
output 	testbus_sel_2;
output 	testbus_sel_3;
input 	sel_enabled_and_granted_1;
input 	pif_enabled_and_granted_1;
output 	reg_plock1;
input 	mutex_grant3;
input 	mutex_grant4;
output 	lif_waitrequest1;
input 	master_read;
input 	wbasic_read_82;
output 	lif_waitrequest2;
output 	basic_reconfig_waitrequest2;
input 	wbasic_writedata_1_8;
input 	wbasic_writedata_2_8;
input 	wbasic_writedata_0_8;
input 	wbasic_writedata_3_8;
output 	lif_number_0;
output 	lif_number_4;
output 	lif_number_3;
output 	lif_number_2;
output 	lif_number_1;
input 	wbasic_writedata_4_8;
input 	wbasic_writedata_5_8;
input 	wbasic_writedata_6_8;
input 	wbasic_writedata_7_8;
input 	wbasic_writedata_8_8;
input 	wbasic_writedata_9_8;
input 	wbasic_writedata_10_8;
input 	wbasic_writedata_11_8;
input 	master_writedata_121;
input 	master_write_data_12;
input 	master_writedata_122;
input 	master_writedata_131;
input 	master_write_data_13;
input 	master_writedata_132;
input 	master_writedata_141;
input 	master_write_data_14;
input 	master_writedata_142;
input 	master_writedata_151;
input 	master_write_data_15;
input 	master_writedata_152;
input 	wbasic_write_83;
input 	lif_is_active;
input 	GND_port;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_from_xcvr_0;
input 	reconfig_from_xcvr_46;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_from_xcvr_1;
input 	reconfig_from_xcvr_47;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_from_xcvr_2;
input 	reconfig_from_xcvr_48;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_from_xcvr_3;
input 	reconfig_from_xcvr_49;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_from_xcvr_4;
input 	reconfig_from_xcvr_50;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_from_xcvr_5;
input 	reconfig_from_xcvr_51;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_from_xcvr_6;
input 	reconfig_from_xcvr_52;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_from_xcvr_7;
input 	reconfig_from_xcvr_53;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_from_xcvr_8;
input 	reconfig_from_xcvr_54;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_from_xcvr_9;
input 	reconfig_from_xcvr_55;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_from_xcvr_10;
input 	reconfig_from_xcvr_56;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_from_xcvr_11;
input 	reconfig_from_xcvr_57;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_from_xcvr_12;
input 	reconfig_from_xcvr_58;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_from_xcvr_13;
input 	reconfig_from_xcvr_59;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_from_xcvr_14;
input 	reconfig_from_xcvr_60;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;
input 	reconfig_from_xcvr_15;
input 	reconfig_from_xcvr_61;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a0~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a1~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a2~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a3~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a16~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a17~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a18~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a19~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a20~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a4~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a21~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a5~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a22~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a6~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a23~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a7~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a24~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a8~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a25~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a9~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a26~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a10~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a27~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a11~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a28~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a12~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a29~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a13~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a30~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a14~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a31~PORTBDATAOUT0 ;
wire \l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a15~PORTBDATAOUT0 ;
wire \l2paddr|physical_addr[11]~q ;
wire \l2paddr|physical_addr[0]~q ;
wire \l2paddr|physical_addr[1]~q ;
wire \l2paddr|physical_addr[2]~q ;
wire \l2paddr|physical_addr[3]~q ;
wire \l2paddr|physical_addr[4]~q ;
wire \l2paddr|physical_addr[5]~q ;
wire \l2paddr|physical_addr[6]~q ;
wire \l2paddr|physical_addr[7]~q ;
wire \l2paddr|physical_addr[8]~q ;
wire \l2paddr|physical_addr[9]~q ;
wire \l2paddr|physical_addr[10]~q ;
wire \Mux19~0_combout ;
wire \Equal12~0_combout ;
wire \always2~0_combout ;
wire \reg_rwdata~0_combout ;
wire \always2~1_combout ;
wire \always2~2_combout ;
wire \reg_rwdata[0]~1_combout ;
wire \reg_rwdata[0]~2_combout ;
wire \reg_rwdata~5_combout ;
wire \reg_rwdata~8_combout ;
wire \reg_rwdata~11_combout ;
wire \reg_rwdata~14_combout ;
wire \reg_rwdata~17_combout ;
wire \reg_rwdata~20_combout ;
wire \reg_rwdata~23_combout ;
wire \reg_rwdata~26_combout ;
wire \reg_rwdata~29_combout ;
wire \reg_rwdata~32_combout ;
wire \reg_rwdata~35_combout ;
wire \reg_rwdata~38_combout ;
wire \reg_rwdata~43_combout ;
wire \reg_rwdata~48_combout ;
wire \reg_rwdata~53_combout ;
wire \always0~0_combout ;
wire \reg_lch[0]~q ;
wire \Mux31~0_combout ;
wire \Add0~1_sumout ;
wire \always1~0_combout ;
wire \lif_inwait~q ;
wire \reg_write_incr~1_combout ;
wire \lif_is_active_last~q ;
wire \reg_write_incr~0_combout ;
wire \reg_write_incr~q ;
wire \reg_addr[2]~0_combout ;
wire \reg_addr[0]~q ;
wire \Mux31~1_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \reg_addr[1]~q ;
wire \reg_lch[1]~q ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \reg_addr[2]~q ;
wire \reg_lch[2]~q ;
wire \reg_is_phys_addr~0_combout ;
wire \reg_is_phys_addr~q ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \reg_addr[3]~q ;
wire \reg_lch[3]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \reg_addr[4]~q ;
wire \reg_lch[4]~q ;
wire \Mux27~0_combout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \reg_addr[5]~q ;
wire \Mux26~0_combout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \reg_addr[6]~q ;
wire \Mux25~0_combout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \reg_addr[7]~q ;
wire \Mux24~0_combout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \reg_addr[8]~q ;
wire \Mux23~0_combout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \reg_addr[9]~q ;
wire \Mux22~0_combout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \reg_addr[10]~q ;
wire \Mux21~0_combout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \reg_addr[11]~q ;
wire \Mux20~0_combout ;
wire \lif_waitrequest~2_combout ;
wire \lif_wrwait~0_combout ;
wire \lif_wrwait~q ;
wire \lif_waitrequest~0_combout ;
wire \always6~0_combout ;
wire \reco_read_length_cntr[2]~0_combout ;
wire \reco_read_length_cntr[2]~1_combout ;
wire \reco_read_length_cntr[1]~2_combout ;
wire \reco_read_length_cntr~3_combout ;
wire \lif_waitrequest~3_combout ;
wire \lif_waitrequest~4_combout ;
wire \always9~0_combout ;
wire \reco_addr_load_cntr[0]~2_combout ;
wire \reco_addr_load_cntr[0]~q ;
wire \reco_addr_load_cntr[1]~0_combout ;
wire \reco_addr_load_cntr[1]~1_combout ;
wire \reco_addr_load_cntr[1]~q ;
wire \Add3~6 ;
wire \Add3~10 ;
wire \Add3~14 ;
wire \Add3~18 ;
wire \Add3~22 ;
wire \Add3~26 ;
wire \Add3~30 ;
wire \Add3~34 ;
wire \Add3~38 ;
wire \Add3~42 ;
wire \Add3~46 ;
wire \Add3~1_sumout ;
wire \reco_addr~0_combout ;
wire \reco_addr[11]~1_combout ;
wire \always2~3_combout ;
wire \reg_rwdata~3_combout ;
wire \reg_rwdata~4_combout ;
wire \reg_rwdata~6_combout ;
wire \reg_rwdata~7_combout ;
wire \reg_rwdata~9_combout ;
wire \reg_rwdata~10_combout ;
wire \reg_rwdata~12_combout ;
wire \reg_rwdata~13_combout ;
wire \reg_rwdata~15_combout ;
wire \reg_rwdata~16_combout ;
wire \reg_rwdata~18_combout ;
wire \reg_rwdata~19_combout ;
wire \reg_rwdata~21_combout ;
wire \reg_rwdata~22_combout ;
wire \reg_rwdata~24_combout ;
wire \reg_rwdata~25_combout ;
wire \reg_rwdata~27_combout ;
wire \reg_rwdata~28_combout ;
wire \reg_rwdata~30_combout ;
wire \reg_rwdata~31_combout ;
wire \reg_rwdata~33_combout ;
wire \reg_rwdata~34_combout ;
wire \reg_rwdata~36_combout ;
wire \reg_rwdata~37_combout ;
wire \reg_rwdata~39_combout ;
wire \reg_rwdata~40_combout ;
wire \reg_rwdata~41_combout ;
wire \reg_rwdata~42_combout ;
wire \reg_rwdata~44_combout ;
wire \reg_rwdata~45_combout ;
wire \reg_rwdata~46_combout ;
wire \reg_rwdata~47_combout ;
wire \reg_rwdata~49_combout ;
wire \reg_rwdata~50_combout ;
wire \reg_rwdata~51_combout ;
wire \reg_rwdata~52_combout ;
wire \reg_rwdata~54_combout ;
wire \reg_rwdata~55_combout ;
wire \reg_rwdata~56_combout ;
wire \reg_rwdata~57_combout ;
wire \always7~0_combout ;
wire \reco_write~0_combout ;
wire \always10~0_combout ;
wire \always10~1_combout ;
wire \Add3~5_sumout ;
wire \reco_addr~2_combout ;
wire \Add3~9_sumout ;
wire \reco_addr~3_combout ;
wire \Add3~13_sumout ;
wire \reco_addr~4_combout ;
wire \Add3~17_sumout ;
wire \reco_addr~5_combout ;
wire \Add3~21_sumout ;
wire \reco_addr~6_combout ;
wire \Add3~25_sumout ;
wire \reco_addr~7_combout ;
wire \Add3~29_sumout ;
wire \reco_addr~8_combout ;
wire \Add3~33_sumout ;
wire \reco_addr~9_combout ;
wire \Add3~37_sumout ;
wire \reco_addr~10_combout ;
wire \Add3~41_sumout ;
wire \reco_addr~11_combout ;
wire \Add3~45_sumout ;
wire \reco_addr~12_combout ;
wire \always6~1_combout ;
wire \reg_plock~0_combout ;
wire \reg_plock~1_combout ;


RECONFIGURE_IP_av_xrbasic_l2p_addr l2paddr(
	.ram_block1a0(ram_block1a0),
	.reg_addr_0(\reg_addr[0]~q ),
	.reg_addr_1(\reg_addr[1]~q ),
	.ram_block1a1(ram_block1a1),
	.reg_addr_2(\reg_addr[2]~q ),
	.ram_block1a2(ram_block1a2),
	.reg_addr_3(\reg_addr[3]~q ),
	.reg_addr_4(\reg_addr[4]~q ),
	.reg_addr_5(\reg_addr[5]~q ),
	.reg_addr_6(\reg_addr[6]~q ),
	.reg_addr_7(\reg_addr[7]~q ),
	.reg_addr_8(\reg_addr[8]~q ),
	.reg_addr_9(\reg_addr[9]~q ),
	.reg_addr_10(\reg_addr[10]~q ),
	.reg_addr_11(\reg_addr[11]~q ),
	.physical_addr_11(\l2paddr|physical_addr[11]~q ),
	.physical_addr_0(\l2paddr|physical_addr[0]~q ),
	.physical_addr_1(\l2paddr|physical_addr[1]~q ),
	.physical_addr_2(\l2paddr|physical_addr[2]~q ),
	.physical_addr_3(\l2paddr|physical_addr[3]~q ),
	.physical_addr_4(\l2paddr|physical_addr[4]~q ),
	.physical_addr_5(\l2paddr|physical_addr[5]~q ),
	.physical_addr_6(\l2paddr|physical_addr[6]~q ),
	.physical_addr_7(\l2paddr|physical_addr[7]~q ),
	.physical_addr_8(\l2paddr|physical_addr[8]~q ),
	.physical_addr_9(\l2paddr|physical_addr[9]~q ),
	.physical_addr_10(\l2paddr|physical_addr[10]~q ),
	.mgmt_clk_clk(mgmt_clk_clk));

RECONFIGURE_IP_av_xrbasic_l2p_rom l2pch(
	.ram_block1a0(ram_block1a0),
	.ram_block1a01(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a0~PORTBDATAOUT0 ),
	.reg_addr_0(\reg_addr[0]~q ),
	.reg_addr_1(\reg_addr[1]~q ),
	.ram_block1a1(ram_block1a1),
	.ram_block1a11(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a1~PORTBDATAOUT0 ),
	.ram_block1a2(ram_block1a2),
	.ram_block1a21(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a2~PORTBDATAOUT0 ),
	.ram_block1a3(ram_block1a3),
	.ram_block1a31(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a3~PORTBDATAOUT0 ),
	.ram_block1a16(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a16~PORTBDATAOUT0 ),
	.ram_block1a17(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a17~PORTBDATAOUT0 ),
	.ram_block1a18(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a18~PORTBDATAOUT0 ),
	.ram_block1a19(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a19~PORTBDATAOUT0 ),
	.ram_block1a20(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a20~PORTBDATAOUT0 ),
	.ram_block1a4(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a4~PORTBDATAOUT0 ),
	.ram_block1a211(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a21~PORTBDATAOUT0 ),
	.ram_block1a5(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a5~PORTBDATAOUT0 ),
	.ram_block1a22(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a22~PORTBDATAOUT0 ),
	.ram_block1a6(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a6~PORTBDATAOUT0 ),
	.ram_block1a23(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a23~PORTBDATAOUT0 ),
	.ram_block1a7(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a7~PORTBDATAOUT0 ),
	.ram_block1a24(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a24~PORTBDATAOUT0 ),
	.ram_block1a8(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a8~PORTBDATAOUT0 ),
	.ram_block1a25(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a25~PORTBDATAOUT0 ),
	.ram_block1a9(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a9~PORTBDATAOUT0 ),
	.ram_block1a26(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a26~PORTBDATAOUT0 ),
	.ram_block1a10(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a10~PORTBDATAOUT0 ),
	.ram_block1a27(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a27~PORTBDATAOUT0 ),
	.ram_block1a111(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a11~PORTBDATAOUT0 ),
	.ram_block1a28(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a28~PORTBDATAOUT0 ),
	.ram_block1a12(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a12~PORTBDATAOUT0 ),
	.ram_block1a29(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a29~PORTBDATAOUT0 ),
	.ram_block1a13(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a13~PORTBDATAOUT0 ),
	.ram_block1a30(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a30~PORTBDATAOUT0 ),
	.ram_block1a14(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a14~PORTBDATAOUT0 ),
	.ram_block1a311(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a31~PORTBDATAOUT0 ),
	.ram_block1a15(\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a15~PORTBDATAOUT0 ),
	.reg_lch_0(\reg_lch[0]~q ),
	.reg_lch_1(\reg_lch[1]~q ),
	.reg_lch_2(\reg_lch[2]~q ),
	.reg_lch_3(\reg_lch[3]~q ),
	.reg_lch_4(\reg_lch[4]~q ),
	.GND_port(GND_port),
	.mgmt_clk_clk(mgmt_clk_clk));

dffeas \basic_reconfig_readdata[12] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_12),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_12),
	.prn(vcc));
defparam \basic_reconfig_readdata[12] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[12] .power_up = "low";

dffeas \basic_reconfig_readdata[13] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_13),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_13),
	.prn(vcc));
defparam \basic_reconfig_readdata[13] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[13] .power_up = "low";

dffeas \basic_reconfig_readdata[14] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_14),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_14),
	.prn(vcc));
defparam \basic_reconfig_readdata[14] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[14] .power_up = "low";

dffeas \basic_reconfig_readdata[15] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_15),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_15),
	.prn(vcc));
defparam \basic_reconfig_readdata[15] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[15] .power_up = "low";

dffeas \basic_reconfig_readdata[16] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_16),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_16),
	.prn(vcc));
defparam \basic_reconfig_readdata[16] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[16] .power_up = "low";

dffeas \basic_reconfig_readdata[17] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_17),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_17),
	.prn(vcc));
defparam \basic_reconfig_readdata[17] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[17] .power_up = "low";

dffeas \basic_reconfig_readdata[18] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_18),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_18),
	.prn(vcc));
defparam \basic_reconfig_readdata[18] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[18] .power_up = "low";

dffeas \basic_reconfig_readdata[19] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_19),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_19),
	.prn(vcc));
defparam \basic_reconfig_readdata[19] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[19] .power_up = "low";

dffeas \basic_reconfig_readdata[20] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_20),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_20),
	.prn(vcc));
defparam \basic_reconfig_readdata[20] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[20] .power_up = "low";

dffeas \basic_reconfig_readdata[21] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_21),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_21),
	.prn(vcc));
defparam \basic_reconfig_readdata[21] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[21] .power_up = "low";

dffeas \basic_reconfig_readdata[22] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_22),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_22),
	.prn(vcc));
defparam \basic_reconfig_readdata[22] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[22] .power_up = "low";

dffeas \basic_reconfig_readdata[23] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_23),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_23),
	.prn(vcc));
defparam \basic_reconfig_readdata[23] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[23] .power_up = "low";

dffeas \basic_reconfig_readdata[24] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_24),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_24),
	.prn(vcc));
defparam \basic_reconfig_readdata[24] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[24] .power_up = "low";

dffeas \basic_reconfig_readdata[25] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_25),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_25),
	.prn(vcc));
defparam \basic_reconfig_readdata[25] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[25] .power_up = "low";

dffeas \basic_reconfig_readdata[26] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_26),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_26),
	.prn(vcc));
defparam \basic_reconfig_readdata[26] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[26] .power_up = "low";

dffeas \basic_reconfig_readdata[27] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_27),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_27),
	.prn(vcc));
defparam \basic_reconfig_readdata[27] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[27] .power_up = "low";

dffeas \basic_reconfig_readdata[28] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_28),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_28),
	.prn(vcc));
defparam \basic_reconfig_readdata[28] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[28] .power_up = "low";

dffeas \basic_reconfig_readdata[29] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_29),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_29),
	.prn(vcc));
defparam \basic_reconfig_readdata[29] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[29] .power_up = "low";

dffeas \basic_reconfig_readdata[30] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_30),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_30),
	.prn(vcc));
defparam \basic_reconfig_readdata[30] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[30] .power_up = "low";

dffeas \basic_reconfig_readdata[31] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(reg_rwdata_31),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal12~0_combout ),
	.ena(vcc),
	.q(basic_reconfig_readdata_31),
	.prn(vcc));
defparam \basic_reconfig_readdata[31] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[31] .power_up = "low";

dffeas \reg_rwdata[16] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_16),
	.prn(vcc));
defparam \reg_rwdata[16] .is_wysiwyg = "true";
defparam \reg_rwdata[16] .power_up = "low";

dffeas \reg_rwdata[17] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_17),
	.prn(vcc));
defparam \reg_rwdata[17] .is_wysiwyg = "true";
defparam \reg_rwdata[17] .power_up = "low";

dffeas \reg_rwdata[18] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_18),
	.prn(vcc));
defparam \reg_rwdata[18] .is_wysiwyg = "true";
defparam \reg_rwdata[18] .power_up = "low";

dffeas \reg_rwdata[19] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_19),
	.prn(vcc));
defparam \reg_rwdata[19] .is_wysiwyg = "true";
defparam \reg_rwdata[19] .power_up = "low";

dffeas \reg_rwdata[20] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_20),
	.prn(vcc));
defparam \reg_rwdata[20] .is_wysiwyg = "true";
defparam \reg_rwdata[20] .power_up = "low";

dffeas \reg_rwdata[21] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_21),
	.prn(vcc));
defparam \reg_rwdata[21] .is_wysiwyg = "true";
defparam \reg_rwdata[21] .power_up = "low";

dffeas \reg_rwdata[22] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_22),
	.prn(vcc));
defparam \reg_rwdata[22] .is_wysiwyg = "true";
defparam \reg_rwdata[22] .power_up = "low";

dffeas \reg_rwdata[23] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_23),
	.prn(vcc));
defparam \reg_rwdata[23] .is_wysiwyg = "true";
defparam \reg_rwdata[23] .power_up = "low";

dffeas \reg_rwdata[24] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_24),
	.prn(vcc));
defparam \reg_rwdata[24] .is_wysiwyg = "true";
defparam \reg_rwdata[24] .power_up = "low";

dffeas \reg_rwdata[25] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_25),
	.prn(vcc));
defparam \reg_rwdata[25] .is_wysiwyg = "true";
defparam \reg_rwdata[25] .power_up = "low";

dffeas \reg_rwdata[26] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_26),
	.prn(vcc));
defparam \reg_rwdata[26] .is_wysiwyg = "true";
defparam \reg_rwdata[26] .power_up = "low";

dffeas \reg_rwdata[27] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_27),
	.prn(vcc));
defparam \reg_rwdata[27] .is_wysiwyg = "true";
defparam \reg_rwdata[27] .power_up = "low";

dffeas \reg_rwdata[28] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_28),
	.prn(vcc));
defparam \reg_rwdata[28] .is_wysiwyg = "true";
defparam \reg_rwdata[28] .power_up = "low";

dffeas \reg_rwdata[29] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_29),
	.prn(vcc));
defparam \reg_rwdata[29] .is_wysiwyg = "true";
defparam \reg_rwdata[29] .power_up = "low";

dffeas \reg_rwdata[30] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_30),
	.prn(vcc));
defparam \reg_rwdata[30] .is_wysiwyg = "true";
defparam \reg_rwdata[30] .power_up = "low";

dffeas \reg_rwdata[31] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~53_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\reg_rwdata[0]~1_combout ),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_31),
	.prn(vcc));
defparam \reg_rwdata[31] .is_wysiwyg = "true";
defparam \reg_rwdata[31] .power_up = "low";

dffeas \basic_reconfig_readdata[0] (
	.clk(mgmt_clk_clk),
	.d(\Mux31~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_0),
	.prn(vcc));
defparam \basic_reconfig_readdata[0] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[0] .power_up = "low";

dffeas \basic_reconfig_readdata[1] (
	.clk(mgmt_clk_clk),
	.d(\Mux30~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_1),
	.prn(vcc));
defparam \basic_reconfig_readdata[1] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[1] .power_up = "low";

dffeas \basic_reconfig_readdata[2] (
	.clk(mgmt_clk_clk),
	.d(\Mux29~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_2),
	.prn(vcc));
defparam \basic_reconfig_readdata[2] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[2] .power_up = "low";

dffeas \basic_reconfig_readdata[3] (
	.clk(mgmt_clk_clk),
	.d(\Mux28~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_3),
	.prn(vcc));
defparam \basic_reconfig_readdata[3] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[3] .power_up = "low";

dffeas \basic_reconfig_readdata[4] (
	.clk(mgmt_clk_clk),
	.d(\Mux27~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_4),
	.prn(vcc));
defparam \basic_reconfig_readdata[4] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[4] .power_up = "low";

dffeas \basic_reconfig_readdata[5] (
	.clk(mgmt_clk_clk),
	.d(\Mux26~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_5),
	.prn(vcc));
defparam \basic_reconfig_readdata[5] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[5] .power_up = "low";

dffeas \basic_reconfig_readdata[6] (
	.clk(mgmt_clk_clk),
	.d(\Mux25~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_6),
	.prn(vcc));
defparam \basic_reconfig_readdata[6] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[6] .power_up = "low";

dffeas \basic_reconfig_readdata[7] (
	.clk(mgmt_clk_clk),
	.d(\Mux24~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_7),
	.prn(vcc));
defparam \basic_reconfig_readdata[7] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[7] .power_up = "low";

dffeas \basic_reconfig_readdata[8] (
	.clk(mgmt_clk_clk),
	.d(\Mux23~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_8),
	.prn(vcc));
defparam \basic_reconfig_readdata[8] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[8] .power_up = "low";

dffeas \basic_reconfig_readdata[9] (
	.clk(mgmt_clk_clk),
	.d(\Mux22~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_9),
	.prn(vcc));
defparam \basic_reconfig_readdata[9] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[9] .power_up = "low";

dffeas \basic_reconfig_readdata[10] (
	.clk(mgmt_clk_clk),
	.d(\Mux21~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_10),
	.prn(vcc));
defparam \basic_reconfig_readdata[10] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[10] .power_up = "low";

dffeas \basic_reconfig_readdata[11] (
	.clk(mgmt_clk_clk),
	.d(\Mux20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(basic_reconfig_readdata_11),
	.prn(vcc));
defparam \basic_reconfig_readdata[11] .is_wysiwyg = "true";
defparam \basic_reconfig_readdata[11] .power_up = "low";

cyclonev_lcell_comb \lif_waitrequest~1 (
	.dataa(!master_write),
	.datab(!wbasic_write_82),
	.datac(!wbasic_address_2_8),
	.datad(!wbasic_address_0_8),
	.datae(!wbasic_address_1_8),
	.dataf(!\lif_waitrequest~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(lif_waitrequest),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_waitrequest~1 .extended_lut = "off";
defparam \lif_waitrequest~1 .lut_mask = 64'h00000D0000000000;
defparam \lif_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \basic_reconfig_waitrequest~0 (
	.dataa(!Equal2),
	.datab(!reconfig_mgmt_read),
	.datac(!mutex_grant),
	.datad(!\lif_inwait~q ),
	.datae(!wbasic_read_8),
	.dataf(!wbasic_read_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(basic_reconfig_waitrequest),
	.sumout(),
	.cout(),
	.shareout());
defparam \basic_reconfig_waitrequest~0 .extended_lut = "off";
defparam \basic_reconfig_waitrequest~0 .lut_mask = 64'h0100FF00FF00FF00;
defparam \basic_reconfig_waitrequest~0 .shared_arith = "off";

dffeas \reco_read_length_cntr[2] (
	.clk(mgmt_clk_clk),
	.d(\reco_read_length_cntr[2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reco_read_length_cntr_2),
	.prn(vcc));
defparam \reco_read_length_cntr[2] .is_wysiwyg = "true";
defparam \reco_read_length_cntr[2] .power_up = "low";

dffeas \reco_read_length_cntr[1] (
	.clk(mgmt_clk_clk),
	.d(\reco_read_length_cntr[1]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reco_read_length_cntr_1),
	.prn(vcc));
defparam \reco_read_length_cntr[1] .is_wysiwyg = "true";
defparam \reco_read_length_cntr[1] .power_up = "low";

dffeas \reco_read_length_cntr[0] (
	.clk(mgmt_clk_clk),
	.d(\reco_read_length_cntr~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reco_read_length_cntr_0),
	.prn(vcc));
defparam \reco_read_length_cntr[0] .is_wysiwyg = "true";
defparam \reco_read_length_cntr[0] .power_up = "low";

cyclonev_lcell_comb \basic_reconfig_waitrequest~1 (
	.dataa(!\lif_waitrequest~2_combout ),
	.datab(!wbasic_address_2_8),
	.datac(!wbasic_address_0_8),
	.datad(!wbasic_address_1_8),
	.datae(!basic_reconfig_waitrequest),
	.dataf(!\lif_waitrequest~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(basic_reconfig_waitrequest1),
	.sumout(),
	.cout(),
	.shareout());
defparam \basic_reconfig_waitrequest~1 .extended_lut = "off";
defparam \basic_reconfig_waitrequest~1 .lut_mask = 64'hFFFB0000FF3B0000;
defparam \basic_reconfig_waitrequest~1 .shared_arith = "off";

dffeas \reco_addr[11] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_11),
	.prn(vcc));
defparam \reco_addr[11] .is_wysiwyg = "true";
defparam \reco_addr[11] .power_up = "low";

dffeas \reg_rwdata[0] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_0),
	.prn(vcc));
defparam \reg_rwdata[0] .is_wysiwyg = "true";
defparam \reg_rwdata[0] .power_up = "low";

dffeas \reg_rwdata[1] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_1),
	.prn(vcc));
defparam \reg_rwdata[1] .is_wysiwyg = "true";
defparam \reg_rwdata[1] .power_up = "low";

dffeas \reg_rwdata[2] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_2),
	.prn(vcc));
defparam \reg_rwdata[2] .is_wysiwyg = "true";
defparam \reg_rwdata[2] .power_up = "low";

dffeas \reg_rwdata[3] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_3),
	.prn(vcc));
defparam \reg_rwdata[3] .is_wysiwyg = "true";
defparam \reg_rwdata[3] .power_up = "low";

dffeas \reg_rwdata[4] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_4),
	.prn(vcc));
defparam \reg_rwdata[4] .is_wysiwyg = "true";
defparam \reg_rwdata[4] .power_up = "low";

dffeas \reg_rwdata[5] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_5),
	.prn(vcc));
defparam \reg_rwdata[5] .is_wysiwyg = "true";
defparam \reg_rwdata[5] .power_up = "low";

dffeas \reg_rwdata[6] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_6),
	.prn(vcc));
defparam \reg_rwdata[6] .is_wysiwyg = "true";
defparam \reg_rwdata[6] .power_up = "low";

dffeas \reg_rwdata[7] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_7),
	.prn(vcc));
defparam \reg_rwdata[7] .is_wysiwyg = "true";
defparam \reg_rwdata[7] .power_up = "low";

dffeas \reg_rwdata[8] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_8),
	.prn(vcc));
defparam \reg_rwdata[8] .is_wysiwyg = "true";
defparam \reg_rwdata[8] .power_up = "low";

dffeas \reg_rwdata[9] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_9),
	.prn(vcc));
defparam \reg_rwdata[9] .is_wysiwyg = "true";
defparam \reg_rwdata[9] .power_up = "low";

dffeas \reg_rwdata[10] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_10),
	.prn(vcc));
defparam \reg_rwdata[10] .is_wysiwyg = "true";
defparam \reg_rwdata[10] .power_up = "low";

dffeas \reg_rwdata[11] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_11),
	.prn(vcc));
defparam \reg_rwdata[11] .is_wysiwyg = "true";
defparam \reg_rwdata[11] .power_up = "low";

dffeas \reg_rwdata[12] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_12),
	.prn(vcc));
defparam \reg_rwdata[12] .is_wysiwyg = "true";
defparam \reg_rwdata[12] .power_up = "low";

dffeas \reg_rwdata[13] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_13),
	.prn(vcc));
defparam \reg_rwdata[13] .is_wysiwyg = "true";
defparam \reg_rwdata[13] .power_up = "low";

dffeas \reg_rwdata[14] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_14),
	.prn(vcc));
defparam \reg_rwdata[14] .is_wysiwyg = "true";
defparam \reg_rwdata[14] .power_up = "low";

dffeas \reg_rwdata[15] (
	.clk(mgmt_clk_clk),
	.d(\reg_rwdata~57_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_rwdata[0]~2_combout ),
	.q(reg_rwdata_15),
	.prn(vcc));
defparam \reg_rwdata[15] .is_wysiwyg = "true";
defparam \reg_rwdata[15] .power_up = "low";

dffeas reco_write(
	.clk(mgmt_clk_clk),
	.d(\reco_write~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reco_write1),
	.prn(vcc));
defparam reco_write.is_wysiwyg = "true";
defparam reco_write.power_up = "low";

dffeas \reco_addr[0] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_0),
	.prn(vcc));
defparam \reco_addr[0] .is_wysiwyg = "true";
defparam \reco_addr[0] .power_up = "low";

dffeas \reco_addr[1] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_1),
	.prn(vcc));
defparam \reco_addr[1] .is_wysiwyg = "true";
defparam \reco_addr[1] .power_up = "low";

dffeas \reco_addr[2] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_2),
	.prn(vcc));
defparam \reco_addr[2] .is_wysiwyg = "true";
defparam \reco_addr[2] .power_up = "low";

dffeas \reco_addr[3] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_3),
	.prn(vcc));
defparam \reco_addr[3] .is_wysiwyg = "true";
defparam \reco_addr[3] .power_up = "low";

dffeas \reco_addr[4] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_4),
	.prn(vcc));
defparam \reco_addr[4] .is_wysiwyg = "true";
defparam \reco_addr[4] .power_up = "low";

dffeas \reco_addr[5] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_5),
	.prn(vcc));
defparam \reco_addr[5] .is_wysiwyg = "true";
defparam \reco_addr[5] .power_up = "low";

dffeas \reco_addr[6] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_6),
	.prn(vcc));
defparam \reco_addr[6] .is_wysiwyg = "true";
defparam \reco_addr[6] .power_up = "low";

dffeas \reco_addr[7] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_7),
	.prn(vcc));
defparam \reco_addr[7] .is_wysiwyg = "true";
defparam \reco_addr[7] .power_up = "low";

dffeas \reco_addr[8] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_8),
	.prn(vcc));
defparam \reco_addr[8] .is_wysiwyg = "true";
defparam \reco_addr[8] .power_up = "low";

dffeas \reco_addr[9] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_9),
	.prn(vcc));
defparam \reco_addr[9] .is_wysiwyg = "true";
defparam \reco_addr[9] .power_up = "low";

dffeas \reco_addr[10] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reco_addr[11]~1_combout ),
	.q(reco_addr_10),
	.prn(vcc));
defparam \reco_addr[10] .is_wysiwyg = "true";
defparam \reco_addr[10] .power_up = "low";

dffeas \testbus_sel[0] (
	.clk(mgmt_clk_clk),
	.d(reg_rwdata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(testbus_sel_0),
	.prn(vcc));
defparam \testbus_sel[0] .is_wysiwyg = "true";
defparam \testbus_sel[0] .power_up = "low";

dffeas \testbus_sel[1] (
	.clk(mgmt_clk_clk),
	.d(reg_rwdata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(testbus_sel_1),
	.prn(vcc));
defparam \testbus_sel[1] .is_wysiwyg = "true";
defparam \testbus_sel[1] .power_up = "low";

dffeas \testbus_sel[2] (
	.clk(mgmt_clk_clk),
	.d(reg_rwdata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(testbus_sel_2),
	.prn(vcc));
defparam \testbus_sel[2] .is_wysiwyg = "true";
defparam \testbus_sel[2] .power_up = "low";

dffeas \testbus_sel[3] (
	.clk(mgmt_clk_clk),
	.d(reg_rwdata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(testbus_sel_3),
	.prn(vcc));
defparam \testbus_sel[3] .is_wysiwyg = "true";
defparam \testbus_sel[3] .power_up = "low";

dffeas reg_plock(
	.clk(mgmt_clk_clk),
	.d(\reg_plock~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reg_plock1),
	.prn(vcc));
defparam reg_plock.is_wysiwyg = "true";
defparam reg_plock.power_up = "low";

cyclonev_lcell_comb \lif_waitrequest~5 (
	.dataa(!master_write),
	.datab(!\lif_inwait~q ),
	.datac(!wbasic_write_82),
	.datad(!wbasic_address_2_8),
	.datae(!wbasic_address_0_8),
	.dataf(!wbasic_address_1_8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(lif_waitrequest1),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_waitrequest~5 .extended_lut = "off";
defparam \lif_waitrequest~5 .lut_mask = 64'h000000000000C400;
defparam \lif_waitrequest~5 .shared_arith = "off";

cyclonev_lcell_comb \lif_waitrequest~6 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!master_read),
	.datae(!\lif_waitrequest~3_combout ),
	.dataf(!wbasic_read_82),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(lif_waitrequest2),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_waitrequest~6 .extended_lut = "off";
defparam \lif_waitrequest~6 .lut_mask = 64'h0808000000080000;
defparam \lif_waitrequest~6 .shared_arith = "off";

cyclonev_lcell_comb \basic_reconfig_waitrequest~2 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(basic_reconfig_waitrequest2),
	.sumout(),
	.cout(),
	.shareout());
defparam \basic_reconfig_waitrequest~2 .extended_lut = "off";
defparam \basic_reconfig_waitrequest~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \basic_reconfig_waitrequest~2 .shared_arith = "off";

dffeas \lif_number[0] (
	.clk(mgmt_clk_clk),
	.d(\reg_lch[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lif_number_0),
	.prn(vcc));
defparam \lif_number[0] .is_wysiwyg = "true";
defparam \lif_number[0] .power_up = "low";

dffeas \lif_number[4] (
	.clk(mgmt_clk_clk),
	.d(\reg_lch[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lif_number_4),
	.prn(vcc));
defparam \lif_number[4] .is_wysiwyg = "true";
defparam \lif_number[4] .power_up = "low";

dffeas \lif_number[3] (
	.clk(mgmt_clk_clk),
	.d(\reg_lch[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lif_number_3),
	.prn(vcc));
defparam \lif_number[3] .is_wysiwyg = "true";
defparam \lif_number[3] .power_up = "low";

dffeas \lif_number[2] (
	.clk(mgmt_clk_clk),
	.d(\reg_lch[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lif_number_2),
	.prn(vcc));
defparam \lif_number[2] .is_wysiwyg = "true";
defparam \lif_number[2] .power_up = "low";

dffeas \lif_number[1] (
	.clk(mgmt_clk_clk),
	.d(\reg_lch[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(lif_number_1),
	.prn(vcc));
defparam \lif_number[1] .is_wysiwyg = "true";
defparam \lif_number[1] .power_up = "low";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "off";
defparam \Mux19~0 .lut_mask = 64'hA1A1A1A1A1A1A1A1;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal12~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal12~0 .extended_lut = "off";
defparam \Equal12~0 .lut_mask = 64'h0808080808080808;
defparam \Equal12~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!master_write),
	.datab(!wbasic_write_82),
	.datac(!wbasic_address_2_8),
	.datad(!wbasic_address_0_8),
	.datae(!wbasic_address_1_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h0000D0000000D000;
defparam \always2~0 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~0 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a16~PORTBDATAOUT0 ),
	.datad(!\always2~0_combout ),
	.datae(!master_writedata_16),
	.dataf(!reconfig_mgmt_writedata_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~0 .extended_lut = "off";
defparam \reg_rwdata~0 .lut_mask = 64'h0F000F330F550F77;
defparam \reg_rwdata~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~1 (
	.dataa(!master_write),
	.datab(!wbasic_write_82),
	.datac(!wbasic_address_2_8),
	.datad(!wbasic_address_0_8),
	.datae(!wbasic_address_1_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'h0D0000000D000000;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \always2~2 (
	.dataa(!wbasic_writedata_1_8),
	.datab(!wbasic_writedata_2_8),
	.datac(!wbasic_writedata_0_8),
	.datad(!wbasic_writedata_3_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~2 .extended_lut = "off";
defparam \always2~2 .lut_mask = 64'h0004000400040004;
defparam \always2~2 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata[0]~1 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~1_combout ),
	.datac(!\always2~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata[0]~1 .extended_lut = "off";
defparam \reg_rwdata[0]~1 .lut_mask = 64'hA8A8A8A8A8A8A8A8;
defparam \reg_rwdata[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata[0]~2 (
	.dataa(!reco_read_length_cntr_2),
	.datab(!reco_read_length_cntr_1),
	.datac(!reco_read_length_cntr_0),
	.datad(!\always2~0_combout ),
	.datae(!\always2~1_combout ),
	.dataf(!\always2~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata[0]~2 .extended_lut = "off";
defparam \reg_rwdata[0]~2 .lut_mask = 64'h20FF20FF20FFFFFF;
defparam \reg_rwdata[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~5 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a17~PORTBDATAOUT0 ),
	.datae(!master_writedata_17),
	.dataf(!reconfig_mgmt_writedata_17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~5 .extended_lut = "off";
defparam \reg_rwdata~5 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~5 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~8 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a18~PORTBDATAOUT0 ),
	.datae(!master_writedata_18),
	.dataf(!reconfig_mgmt_writedata_18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~8 .extended_lut = "off";
defparam \reg_rwdata~8 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~8 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~11 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a19~PORTBDATAOUT0 ),
	.datae(!master_writedata_19),
	.dataf(!reconfig_mgmt_writedata_19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~11 .extended_lut = "off";
defparam \reg_rwdata~11 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~11 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~14 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a20~PORTBDATAOUT0 ),
	.datae(!master_writedata_20),
	.dataf(!reconfig_mgmt_writedata_20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~14 .extended_lut = "off";
defparam \reg_rwdata~14 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~14 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~17 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a21~PORTBDATAOUT0 ),
	.datae(!master_writedata_21),
	.dataf(!reconfig_mgmt_writedata_21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~17 .extended_lut = "off";
defparam \reg_rwdata~17 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~17 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~20 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a22~PORTBDATAOUT0 ),
	.datae(!master_writedata_22),
	.dataf(!reconfig_mgmt_writedata_22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~20 .extended_lut = "off";
defparam \reg_rwdata~20 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~20 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~23 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a23~PORTBDATAOUT0 ),
	.datae(!master_writedata_23),
	.dataf(!reconfig_mgmt_writedata_23),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~23 .extended_lut = "off";
defparam \reg_rwdata~23 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~23 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~26 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a24~PORTBDATAOUT0 ),
	.datae(!master_writedata_24),
	.dataf(!reconfig_mgmt_writedata_24),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~26 .extended_lut = "off";
defparam \reg_rwdata~26 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~26 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~29 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a25~PORTBDATAOUT0 ),
	.datae(!master_writedata_25),
	.dataf(!reconfig_mgmt_writedata_25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~29 .extended_lut = "off";
defparam \reg_rwdata~29 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~29 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~32 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a26~PORTBDATAOUT0 ),
	.datae(!master_writedata_26),
	.dataf(!reconfig_mgmt_writedata_26),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~32 .extended_lut = "off";
defparam \reg_rwdata~32 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~32 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~35 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a27~PORTBDATAOUT0 ),
	.datae(!master_writedata_27),
	.dataf(!reconfig_mgmt_writedata_27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~35 .extended_lut = "off";
defparam \reg_rwdata~35 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~35 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~38 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a28~PORTBDATAOUT0 ),
	.datae(!master_writedata_28),
	.dataf(!reconfig_mgmt_writedata_28),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~38 .extended_lut = "off";
defparam \reg_rwdata~38 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~38 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~43 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a29~PORTBDATAOUT0 ),
	.datae(!master_writedata_29),
	.dataf(!reconfig_mgmt_writedata_29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~43 .extended_lut = "off";
defparam \reg_rwdata~43 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~43 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~48 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a30~PORTBDATAOUT0 ),
	.datae(!master_writedata_30),
	.dataf(!reconfig_mgmt_writedata_30),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~48 .extended_lut = "off";
defparam \reg_rwdata~48 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~48 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~53 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant2),
	.datac(!\always2~0_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a31~PORTBDATAOUT0 ),
	.datae(!master_writedata_31),
	.dataf(!reconfig_mgmt_writedata_31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~53 .extended_lut = "off";
defparam \reg_rwdata~53 .lut_mask = 64'h00F003F305F507F7;
defparam \reg_rwdata~53 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!master_write),
	.datab(!wbasic_write_82),
	.datac(!wbasic_address_2_8),
	.datad(!wbasic_address_0_8),
	.datae(!wbasic_address_1_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h00000D0000000D00;
defparam \always0~0 .shared_arith = "off";

dffeas \reg_lch[0] (
	.clk(mgmt_clk_clk),
	.d(wbasic_writedata_0_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\reg_lch[0]~q ),
	.prn(vcc));
defparam \reg_lch[0] .is_wysiwyg = "true";
defparam \reg_lch[0] .power_up = "low";

cyclonev_lcell_comb \Mux31~0 (
	.dataa(!wbasic_address_0_8),
	.datab(!wbasic_address_1_8),
	.datac(!pif_enabled_and_granted_0),
	.datad(!pif_enabled_and_granted_1),
	.datae(!ram_block1a0),
	.dataf(!\reg_lch[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~0 .extended_lut = "off";
defparam \Mux31~0 .lut_mask = 64'hE666A222C4448000;
defparam \Mux31~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!wbasic_write_83),
	.datab(!wbasic_address_2_8),
	.datac(!wbasic_address_0_8),
	.datad(!wbasic_address_1_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'h0008000800080008;
defparam \always1~0 .shared_arith = "off";

dffeas lif_inwait(
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_waitrequest2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lif_inwait~q ),
	.prn(vcc));
defparam lif_inwait.is_wysiwyg = "true";
defparam lif_inwait.power_up = "low";

cyclonev_lcell_comb \reg_write_incr~1 (
	.dataa(!\reg_write_incr~q ),
	.datab(!wbasic_writedata_1_8),
	.datac(!wbasic_writedata_2_8),
	.datad(!wbasic_writedata_0_8),
	.datae(!wbasic_writedata_3_8),
	.dataf(!\always2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_write_incr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_write_incr~1 .extended_lut = "off";
defparam \reg_write_incr~1 .lut_mask = 64'h0000000054575555;
defparam \reg_write_incr~1 .shared_arith = "off";

dffeas lif_is_active_last(
	.clk(mgmt_clk_clk),
	.d(lif_is_active),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lif_is_active_last~q ),
	.prn(vcc));
defparam lif_is_active_last.is_wysiwyg = "true";
defparam lif_is_active_last.power_up = "low";

cyclonev_lcell_comb \reg_write_incr~0 (
	.dataa(!\always2~1_combout ),
	.datab(!\lif_is_active_last~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_write_incr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_write_incr~0 .extended_lut = "off";
defparam \reg_write_incr~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \reg_write_incr~0 .shared_arith = "off";

dffeas reg_write_incr(
	.clk(mgmt_clk_clk),
	.d(\reg_write_incr~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_write_incr~0_combout ),
	.q(\reg_write_incr~q ),
	.prn(vcc));
defparam reg_write_incr.is_wysiwyg = "true";
defparam reg_write_incr.power_up = "low";

cyclonev_lcell_comb \reg_addr[2]~0 (
	.dataa(!\lif_inwait~q ),
	.datab(!wbasic_write_83),
	.datac(!wbasic_address_2_8),
	.datad(!wbasic_address_0_8),
	.datae(!wbasic_address_1_8),
	.dataf(!\reg_write_incr~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_addr[2]~0 .extended_lut = "off";
defparam \reg_addr[2]~0 .lut_mask = 64'h000000C0000080C0;
defparam \reg_addr[2]~0 .shared_arith = "off";

dffeas \reg_addr[0] (
	.clk(mgmt_clk_clk),
	.d(\Add0~1_sumout ),
	.asdata(wbasic_writedata_0_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[0]~q ),
	.prn(vcc));
defparam \reg_addr[0] .is_wysiwyg = "true";
defparam \reg_addr[0] .power_up = "low";

cyclonev_lcell_comb \Mux31~1 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_0),
	.datae(!\Mux31~0_combout ),
	.dataf(!\reg_addr[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux31~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~1 .extended_lut = "off";
defparam \Mux31~1 .lut_mask = 64'hF5FDA0A8F7FFA2AA;
defparam \Mux31~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \reg_addr[1] (
	.clk(mgmt_clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(wbasic_writedata_1_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[1]~q ),
	.prn(vcc));
defparam \reg_addr[1] .is_wysiwyg = "true";
defparam \reg_addr[1] .power_up = "low";

dffeas \reg_lch[1] (
	.clk(mgmt_clk_clk),
	.d(wbasic_writedata_1_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\reg_lch[1]~q ),
	.prn(vcc));
defparam \reg_lch[1] .is_wysiwyg = "true";
defparam \reg_lch[1] .power_up = "low";

cyclonev_lcell_comb \Mux30~0 (
	.dataa(!wbasic_address_0_8),
	.datab(!wbasic_address_1_8),
	.datac(!ram_block1a1),
	.datad(!\reg_lch[1]~q ),
	.datae(!reg_plock1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~0 .extended_lut = "off";
defparam \Mux30~0 .lut_mask = 64'hEAC86240EAC86240;
defparam \Mux30~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux30~1 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_1),
	.datae(!\reg_addr[1]~q ),
	.dataf(!\Mux30~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux30~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~1 .extended_lut = "off";
defparam \Mux30~1 .lut_mask = 64'hF5FDF7FFA0A8A2AA;
defparam \Mux30~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \reg_addr[2] (
	.clk(mgmt_clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(wbasic_writedata_2_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[2]~q ),
	.prn(vcc));
defparam \reg_addr[2] .is_wysiwyg = "true";
defparam \reg_addr[2] .power_up = "low";

dffeas \reg_lch[2] (
	.clk(mgmt_clk_clk),
	.d(wbasic_writedata_2_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\reg_lch[2]~q ),
	.prn(vcc));
defparam \reg_lch[2] .is_wysiwyg = "true";
defparam \reg_lch[2] .power_up = "low";

cyclonev_lcell_comb \reg_is_phys_addr~0 (
	.dataa(!\reg_is_phys_addr~q ),
	.datab(!wbasic_writedata_1_8),
	.datac(!wbasic_writedata_2_8),
	.datad(!wbasic_writedata_0_8),
	.datae(!wbasic_writedata_3_8),
	.dataf(!\always2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_is_phys_addr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_is_phys_addr~0 .extended_lut = "off";
defparam \reg_is_phys_addr~0 .lut_mask = 64'h0000000045755555;
defparam \reg_is_phys_addr~0 .shared_arith = "off";

dffeas reg_is_phys_addr(
	.clk(mgmt_clk_clk),
	.d(\reg_is_phys_addr~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reg_write_incr~0_combout ),
	.q(\reg_is_phys_addr~q ),
	.prn(vcc));
defparam reg_is_phys_addr.is_wysiwyg = "true";
defparam reg_is_phys_addr.power_up = "low";

cyclonev_lcell_comb \Mux29~0 (
	.dataa(!wbasic_address_0_8),
	.datab(!wbasic_address_1_8),
	.datac(!ram_block1a2),
	.datad(!\reg_lch[2]~q ),
	.datae(!\reg_is_phys_addr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~0 .extended_lut = "off";
defparam \Mux29~0 .lut_mask = 64'hEAC86240EAC86240;
defparam \Mux29~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux29~1 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_2),
	.datae(!\reg_addr[2]~q ),
	.dataf(!\Mux29~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux29~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~1 .extended_lut = "off";
defparam \Mux29~1 .lut_mask = 64'hF5FDF7FFA0A8A2AA;
defparam \Mux29~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \reg_addr[3] (
	.clk(mgmt_clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(wbasic_writedata_3_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[3]~q ),
	.prn(vcc));
defparam \reg_addr[3] .is_wysiwyg = "true";
defparam \reg_addr[3] .power_up = "low";

dffeas \reg_lch[3] (
	.clk(mgmt_clk_clk),
	.d(wbasic_writedata_3_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\reg_lch[3]~q ),
	.prn(vcc));
defparam \reg_lch[3] .is_wysiwyg = "true";
defparam \reg_lch[3] .power_up = "low";

cyclonev_lcell_comb \Mux28~0 (
	.dataa(!wbasic_address_0_8),
	.datab(!wbasic_address_1_8),
	.datac(!ram_block1a3),
	.datad(!\reg_lch[3]~q ),
	.datae(!\reg_write_incr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~0 .extended_lut = "off";
defparam \Mux28~0 .lut_mask = 64'hEAC86240EAC86240;
defparam \Mux28~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~1 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_3),
	.datae(!\reg_addr[3]~q ),
	.dataf(!\Mux28~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~1 .extended_lut = "off";
defparam \Mux28~1 .lut_mask = 64'hF5FDF7FFA0A8A2AA;
defparam \Mux28~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \reg_addr[4] (
	.clk(mgmt_clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(wbasic_writedata_4_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[4]~q ),
	.prn(vcc));
defparam \reg_addr[4] .is_wysiwyg = "true";
defparam \reg_addr[4] .power_up = "low";

dffeas \reg_lch[4] (
	.clk(mgmt_clk_clk),
	.d(wbasic_writedata_4_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\reg_lch[4]~q ),
	.prn(vcc));
defparam \reg_lch[4] .is_wysiwyg = "true";
defparam \reg_lch[4] .power_up = "low";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_4),
	.datae(!\reg_addr[4]~q ),
	.dataf(!\reg_lch[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "off";
defparam \Mux27~0 .lut_mask = 64'hA1A9A3ABA5ADA7AF;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \reg_addr[5] (
	.clk(mgmt_clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(wbasic_writedata_5_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[5]~q ),
	.prn(vcc));
defparam \reg_addr[5] .is_wysiwyg = "true";
defparam \reg_addr[5] .power_up = "low";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_5),
	.datae(!\reg_addr[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "off";
defparam \Mux26~0 .lut_mask = 64'hA1A9A3ABA1A9A3AB;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \reg_addr[6] (
	.clk(mgmt_clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(wbasic_writedata_6_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[6]~q ),
	.prn(vcc));
defparam \reg_addr[6] .is_wysiwyg = "true";
defparam \reg_addr[6] .power_up = "low";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_6),
	.datae(!\reg_addr[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "off";
defparam \Mux25~0 .lut_mask = 64'hA1A9A3ABA1A9A3AB;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \reg_addr[7] (
	.clk(mgmt_clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(wbasic_writedata_7_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[7]~q ),
	.prn(vcc));
defparam \reg_addr[7] .is_wysiwyg = "true";
defparam \reg_addr[7] .power_up = "low";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_7),
	.datae(!\reg_addr[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "off";
defparam \Mux24~0 .lut_mask = 64'hA1A9A3ABA1A9A3AB;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \reg_addr[8] (
	.clk(mgmt_clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(wbasic_writedata_8_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[8]~q ),
	.prn(vcc));
defparam \reg_addr[8] .is_wysiwyg = "true";
defparam \reg_addr[8] .power_up = "low";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_8),
	.datae(!\reg_addr[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "off";
defparam \Mux23~0 .lut_mask = 64'hA1A9A3ABA1A9A3AB;
defparam \Mux23~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \reg_addr[9] (
	.clk(mgmt_clk_clk),
	.d(\Add0~37_sumout ),
	.asdata(wbasic_writedata_9_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[9]~q ),
	.prn(vcc));
defparam \reg_addr[9] .is_wysiwyg = "true";
defparam \reg_addr[9] .power_up = "low";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_9),
	.datae(!\reg_addr[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "off";
defparam \Mux22~0 .lut_mask = 64'hA1A9A3ABA1A9A3AB;
defparam \Mux22~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \reg_addr[10] (
	.clk(mgmt_clk_clk),
	.d(\Add0~41_sumout ),
	.asdata(wbasic_writedata_10_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[10]~q ),
	.prn(vcc));
defparam \reg_addr[10] .is_wysiwyg = "true";
defparam \reg_addr[10] .power_up = "low";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_10),
	.datae(!\reg_addr[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "off";
defparam \Mux21~0 .lut_mask = 64'hA1A9A3ABA1A9A3AB;
defparam \Mux21~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\reg_addr[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \reg_addr[11] (
	.clk(mgmt_clk_clk),
	.d(\Add0~45_sumout ),
	.asdata(wbasic_writedata_11_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always1~0_combout ),
	.ena(\reg_addr[2]~0_combout ),
	.q(\reg_addr[11]~q ),
	.prn(vcc));
defparam \reg_addr[11] .is_wysiwyg = "true";
defparam \reg_addr[11] .power_up = "low";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(!reg_rwdata_11),
	.datae(!\reg_addr[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "off";
defparam \Mux20~0 .lut_mask = 64'hA1A9A3ABA1A9A3AB;
defparam \Mux20~0 .shared_arith = "off";

cyclonev_lcell_comb \lif_waitrequest~2 (
	.dataa(!Equal2),
	.datab(!mutex_grant),
	.datac(!reconfig_mgmt_write),
	.datad(!\lif_inwait~q ),
	.datae(!wbasic_write_8),
	.dataf(!wbasic_write_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_waitrequest~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_waitrequest~2 .extended_lut = "off";
defparam \lif_waitrequest~2 .lut_mask = 64'h0100FF00FF00FF00;
defparam \lif_waitrequest~2 .shared_arith = "off";

cyclonev_lcell_comb \lif_wrwait~0 (
	.dataa(!\lif_waitrequest~2_combout ),
	.datab(!wbasic_address_2_8),
	.datac(!wbasic_address_0_8),
	.datad(!wbasic_address_1_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_wrwait~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_wrwait~0 .extended_lut = "off";
defparam \lif_wrwait~0 .lut_mask = 64'h0010001000100010;
defparam \lif_wrwait~0 .shared_arith = "off";

dffeas lif_wrwait(
	.clk(mgmt_clk_clk),
	.d(\lif_wrwait~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lif_wrwait~q ),
	.prn(vcc));
defparam lif_wrwait.is_wysiwyg = "true";
defparam lif_wrwait.power_up = "low";

cyclonev_lcell_comb \lif_waitrequest~0 (
	.dataa(!\lif_inwait~q ),
	.datab(!\lif_wrwait~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_waitrequest~0 .extended_lut = "off";
defparam \lif_waitrequest~0 .lut_mask = 64'h4444444444444444;
defparam \lif_waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \always6~0 (
	.dataa(!\lif_waitrequest~2_combout ),
	.datab(!wbasic_address_2_8),
	.datac(!wbasic_address_0_8),
	.datad(!wbasic_address_1_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'h1000100010001000;
defparam \always6~0 .shared_arith = "off";

cyclonev_lcell_comb \reco_read_length_cntr[2]~0 (
	.dataa(!\always6~0_combout ),
	.datab(!wbasic_writedata_1_8),
	.datac(!wbasic_writedata_2_8),
	.datad(!wbasic_writedata_0_8),
	.datae(!wbasic_writedata_3_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_read_length_cntr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_read_length_cntr[2]~0 .extended_lut = "off";
defparam \reco_read_length_cntr[2]~0 .lut_mask = 64'h0040000000400000;
defparam \reco_read_length_cntr[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \reco_read_length_cntr[2]~1 (
	.dataa(!reco_read_length_cntr_2),
	.datab(!reco_read_length_cntr_1),
	.datac(!reco_read_length_cntr_0),
	.datad(!\reco_read_length_cntr[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_read_length_cntr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_read_length_cntr[2]~1 .extended_lut = "off";
defparam \reco_read_length_cntr[2]~1 .lut_mask = 64'h15FF15FF15FF15FF;
defparam \reco_read_length_cntr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \reco_read_length_cntr[1]~2 (
	.dataa(!reco_read_length_cntr_2),
	.datab(!reco_read_length_cntr_1),
	.datac(!reco_read_length_cntr_0),
	.datad(!\reco_read_length_cntr[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_read_length_cntr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_read_length_cntr[1]~2 .extended_lut = "off";
defparam \reco_read_length_cntr[1]~2 .lut_mask = 64'h43FF43FF43FF43FF;
defparam \reco_read_length_cntr[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \reco_read_length_cntr~3 (
	.dataa(!reco_read_length_cntr_2),
	.datab(!reco_read_length_cntr_1),
	.datac(!reco_read_length_cntr_0),
	.datad(!\reco_read_length_cntr[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_read_length_cntr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_read_length_cntr~3 .extended_lut = "off";
defparam \reco_read_length_cntr~3 .lut_mask = 64'h7000700070007000;
defparam \reco_read_length_cntr~3 .shared_arith = "off";

cyclonev_lcell_comb \lif_waitrequest~3 (
	.dataa(!reco_read_length_cntr_2),
	.datab(!reco_read_length_cntr_1),
	.datac(!reco_read_length_cntr_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_waitrequest~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_waitrequest~3 .extended_lut = "off";
defparam \lif_waitrequest~3 .lut_mask = 64'h8080808080808080;
defparam \lif_waitrequest~3 .shared_arith = "off";

cyclonev_lcell_comb \lif_waitrequest~4 (
	.dataa(!Equal2),
	.datab(!reconfig_mgmt_read),
	.datac(!mutex_grant),
	.datad(!\lif_waitrequest~3_combout ),
	.datae(!wbasic_read_8),
	.dataf(!wbasic_read_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lif_waitrequest~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lif_waitrequest~4 .extended_lut = "off";
defparam \lif_waitrequest~4 .lut_mask = 64'h0100FF00FF00FF00;
defparam \lif_waitrequest~4 .shared_arith = "off";

cyclonev_lcell_comb \always9~0 (
	.dataa(!\always6~0_combout ),
	.datab(!wbasic_writedata_1_8),
	.datac(!wbasic_writedata_2_8),
	.datad(!wbasic_writedata_3_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~0 .extended_lut = "off";
defparam \always9~0 .lut_mask = 64'h1000100010001000;
defparam \always9~0 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr_load_cntr[0]~2 (
	.dataa(!lif_waitrequest1),
	.datab(!\lif_wrwait~0_combout ),
	.datac(!\reco_addr_load_cntr[1]~q ),
	.datad(!\reco_addr_load_cntr[0]~q ),
	.datae(!\always9~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr_load_cntr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr_load_cntr[0]~2 .extended_lut = "off";
defparam \reco_addr_load_cntr[0]~2 .lut_mask = 64'h3B33BBBB3B33BBBB;
defparam \reco_addr_load_cntr[0]~2 .shared_arith = "off";

dffeas \reco_addr_load_cntr[0] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr_load_cntr[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reco_addr_load_cntr[0]~q ),
	.prn(vcc));
defparam \reco_addr_load_cntr[0] .is_wysiwyg = "true";
defparam \reco_addr_load_cntr[0] .power_up = "low";

cyclonev_lcell_comb \reco_addr_load_cntr[1]~0 (
	.dataa(!wbasic_address_2_8),
	.datab(!wbasic_address_0_8),
	.datac(!wbasic_address_1_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr_load_cntr[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr_load_cntr[1]~0 .extended_lut = "off";
defparam \reco_addr_load_cntr[1]~0 .lut_mask = 64'h0606060606060606;
defparam \reco_addr_load_cntr[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr_load_cntr[1]~1 (
	.dataa(!\lif_waitrequest~2_combout ),
	.datab(!\reco_addr_load_cntr[1]~q ),
	.datac(!\reco_addr_load_cntr[0]~q ),
	.datad(!\always9~0_combout ),
	.datae(!\reco_addr_load_cntr[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr_load_cntr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr_load_cntr[1]~1 .extended_lut = "off";
defparam \reco_addr_load_cntr[1]~1 .lut_mask = 64'h0302575703025757;
defparam \reco_addr_load_cntr[1]~1 .shared_arith = "off";

dffeas \reco_addr_load_cntr[1] (
	.clk(mgmt_clk_clk),
	.d(\reco_addr_load_cntr[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reco_addr_load_cntr[1]~q ),
	.prn(vcc));
defparam \reco_addr_load_cntr[1] .is_wysiwyg = "true";
defparam \reco_addr_load_cntr[1] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h00000000000000FF;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~9 .shared_arith = "off";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~13 .shared_arith = "off";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~17 .shared_arith = "off";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~21 .shared_arith = "off";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~25 .shared_arith = "off";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~29 .shared_arith = "off";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~33 .shared_arith = "off";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout());
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~37 .shared_arith = "off";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout());
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~41 .shared_arith = "off";

cyclonev_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout());
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~45 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reco_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~0 (
	.dataa(!\reg_is_phys_addr~q ),
	.datab(!\reg_addr[11]~q ),
	.datac(!\l2paddr|physical_addr[11]~q ),
	.datad(!\reco_addr_load_cntr[1]~q ),
	.datae(!\reco_addr_load_cntr[0]~q ),
	.dataf(!\Add3~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~0 .extended_lut = "off";
defparam \reco_addr~0 .lut_mask = 64'h00003B00FFFF3BFF;
defparam \reco_addr~0 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr[11]~1 (
	.dataa(!reco_write1),
	.datab(!\reg_write_incr~q ),
	.datac(!\reco_addr_load_cntr[1]~q ),
	.datad(!\reco_addr_load_cntr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr[11]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr[11]~1 .extended_lut = "off";
defparam \reco_addr[11]~1 .lut_mask = 64'h11F111F111F111F1;
defparam \reco_addr[11]~1 .shared_arith = "off";

cyclonev_lcell_comb \always2~3 (
	.dataa(!\always2~1_combout ),
	.datab(!\always2~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~3 .extended_lut = "off";
defparam \always2~3 .lut_mask = 64'h1111111111111111;
defparam \always2~3 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~3 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_0),
	.datad(!reconfig_from_xcvr_46),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~3 .extended_lut = "off";
defparam \reg_rwdata~3 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~3 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~4 (
	.dataa(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a0~PORTBDATAOUT0 ),
	.datab(!wbasic_writedata_0_8),
	.datac(!\always2~0_combout ),
	.datad(!\always2~3_combout ),
	.datae(!\reg_rwdata~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~4 .extended_lut = "off";
defparam \reg_rwdata~4 .lut_mask = 64'h0353F3530353F353;
defparam \reg_rwdata~4 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~6 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_1),
	.datad(!reconfig_from_xcvr_47),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~6 .extended_lut = "off";
defparam \reg_rwdata~6 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~6 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~7 (
	.dataa(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a1~PORTBDATAOUT0 ),
	.datab(!wbasic_writedata_1_8),
	.datac(!\always2~0_combout ),
	.datad(!\always2~3_combout ),
	.datae(!\reg_rwdata~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~7 .extended_lut = "off";
defparam \reg_rwdata~7 .lut_mask = 64'h0353F3530353F353;
defparam \reg_rwdata~7 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~9 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_2),
	.datad(!reconfig_from_xcvr_48),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~9 .extended_lut = "off";
defparam \reg_rwdata~9 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~9 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~10 (
	.dataa(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a2~PORTBDATAOUT0 ),
	.datab(!wbasic_writedata_2_8),
	.datac(!\always2~0_combout ),
	.datad(!\always2~3_combout ),
	.datae(!\reg_rwdata~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~10 .extended_lut = "off";
defparam \reg_rwdata~10 .lut_mask = 64'h0353F3530353F353;
defparam \reg_rwdata~10 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~12 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_3),
	.datad(!reconfig_from_xcvr_49),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~12 .extended_lut = "off";
defparam \reg_rwdata~12 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~12 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~13 (
	.dataa(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a3~PORTBDATAOUT0 ),
	.datab(!wbasic_writedata_3_8),
	.datac(!\always2~0_combout ),
	.datad(!\always2~3_combout ),
	.datae(!\reg_rwdata~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~13 .extended_lut = "off";
defparam \reg_rwdata~13 .lut_mask = 64'h0353F3530353F353;
defparam \reg_rwdata~13 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~15 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_4),
	.datad(!reconfig_from_xcvr_50),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~15 .extended_lut = "off";
defparam \reg_rwdata~15 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~15 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~16 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_4_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a4~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~16 .extended_lut = "off";
defparam \reg_rwdata~16 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~16 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~18 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_5),
	.datad(!reconfig_from_xcvr_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~18 .extended_lut = "off";
defparam \reg_rwdata~18 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~18 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~19 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_5_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a5~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~19 .extended_lut = "off";
defparam \reg_rwdata~19 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~19 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~21 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_6),
	.datad(!reconfig_from_xcvr_52),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~21 .extended_lut = "off";
defparam \reg_rwdata~21 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~21 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~22 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_6_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a6~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~22 .extended_lut = "off";
defparam \reg_rwdata~22 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~22 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~24 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_7),
	.datad(!reconfig_from_xcvr_53),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~24 .extended_lut = "off";
defparam \reg_rwdata~24 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~24 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~25 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_7_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a7~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~25 .extended_lut = "off";
defparam \reg_rwdata~25 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~25 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~27 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_8),
	.datad(!reconfig_from_xcvr_54),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~27 .extended_lut = "off";
defparam \reg_rwdata~27 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~27 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~28 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_8_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a8~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~28 .extended_lut = "off";
defparam \reg_rwdata~28 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~28 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~30 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_9),
	.datad(!reconfig_from_xcvr_55),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~30 .extended_lut = "off";
defparam \reg_rwdata~30 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~30 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~31 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_9_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a9~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~31 .extended_lut = "off";
defparam \reg_rwdata~31 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~31 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~33 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_10),
	.datad(!reconfig_from_xcvr_56),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~33 .extended_lut = "off";
defparam \reg_rwdata~33 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~33 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~34 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_10_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a10~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~34 .extended_lut = "off";
defparam \reg_rwdata~34 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~34 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~36 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!reconfig_from_xcvr_11),
	.datad(!reconfig_from_xcvr_57),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~36 .extended_lut = "off";
defparam \reg_rwdata~36 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~36 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~37 (
	.dataa(!\always2~0_combout ),
	.datab(!\always2~3_combout ),
	.datac(!wbasic_writedata_11_8),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a11~PORTBDATAOUT0 ),
	.datae(!\reg_rwdata~36_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~37 .extended_lut = "off";
defparam \reg_rwdata~37 .lut_mask = 64'h05278DAF05278DAF;
defparam \reg_rwdata~37 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~39 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant1),
	.datac(!reconfig_mgmt_writedata_12),
	.datad(!master_writedata_122),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~39 .extended_lut = "off";
defparam \reg_rwdata~39 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~39 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~40 (
	.dataa(!mutex_grant4),
	.datab(!mutex_grant2),
	.datac(!master_write_data_12),
	.datad(!master_writedata_12),
	.datae(!\reg_rwdata~39_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~40 .extended_lut = "off";
defparam \reg_rwdata~40 .lut_mask = 64'hFAC80000FAC80000;
defparam \reg_rwdata~40 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~41 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!\always2~3_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a12~PORTBDATAOUT0 ),
	.datae(!reconfig_from_xcvr_12),
	.dataf(!reconfig_from_xcvr_58),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~41 .extended_lut = "off";
defparam \reg_rwdata~41 .lut_mask = 64'h000F505F303F707F;
defparam \reg_rwdata~41 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~42 (
	.dataa(!mutex_grant3),
	.datab(!\always2~0_combout ),
	.datac(!master_writedata_121),
	.datad(!\reg_rwdata~40_combout ),
	.datae(!\reg_rwdata~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~42 .extended_lut = "off";
defparam \reg_rwdata~42 .lut_mask = 64'h3301FFCD3301FFCD;
defparam \reg_rwdata~42 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~44 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant1),
	.datac(!reconfig_mgmt_writedata_13),
	.datad(!master_writedata_132),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~44 .extended_lut = "off";
defparam \reg_rwdata~44 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~44 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~45 (
	.dataa(!mutex_grant4),
	.datab(!mutex_grant2),
	.datac(!master_write_data_13),
	.datad(!master_writedata_13),
	.datae(!\reg_rwdata~44_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~45 .extended_lut = "off";
defparam \reg_rwdata~45 .lut_mask = 64'hFAC80000FAC80000;
defparam \reg_rwdata~45 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~46 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!\always2~3_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a13~PORTBDATAOUT0 ),
	.datae(!reconfig_from_xcvr_13),
	.dataf(!reconfig_from_xcvr_59),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~46 .extended_lut = "off";
defparam \reg_rwdata~46 .lut_mask = 64'h000F505F303F707F;
defparam \reg_rwdata~46 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~47 (
	.dataa(!mutex_grant3),
	.datab(!\always2~0_combout ),
	.datac(!master_writedata_131),
	.datad(!\reg_rwdata~45_combout ),
	.datae(!\reg_rwdata~46_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~47 .extended_lut = "off";
defparam \reg_rwdata~47 .lut_mask = 64'h3301FFCD3301FFCD;
defparam \reg_rwdata~47 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~49 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant1),
	.datac(!reconfig_mgmt_writedata_14),
	.datad(!master_writedata_142),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~49 .extended_lut = "off";
defparam \reg_rwdata~49 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~49 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~50 (
	.dataa(!mutex_grant4),
	.datab(!mutex_grant2),
	.datac(!master_write_data_14),
	.datad(!master_writedata_14),
	.datae(!\reg_rwdata~49_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~50 .extended_lut = "off";
defparam \reg_rwdata~50 .lut_mask = 64'hFAC80000FAC80000;
defparam \reg_rwdata~50 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~51 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!\always2~3_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a14~PORTBDATAOUT0 ),
	.datae(!reconfig_from_xcvr_14),
	.dataf(!reconfig_from_xcvr_60),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~51 .extended_lut = "off";
defparam \reg_rwdata~51 .lut_mask = 64'h000F505F303F707F;
defparam \reg_rwdata~51 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~52 (
	.dataa(!mutex_grant3),
	.datab(!\always2~0_combout ),
	.datac(!master_writedata_141),
	.datad(!\reg_rwdata~50_combout ),
	.datae(!\reg_rwdata~51_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~52 .extended_lut = "off";
defparam \reg_rwdata~52 .lut_mask = 64'h3301FFCD3301FFCD;
defparam \reg_rwdata~52 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~54 (
	.dataa(!mutex_grant),
	.datab(!mutex_grant1),
	.datac(!reconfig_mgmt_writedata_15),
	.datad(!master_writedata_152),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~54 .extended_lut = "off";
defparam \reg_rwdata~54 .lut_mask = 64'h0537053705370537;
defparam \reg_rwdata~54 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~55 (
	.dataa(!mutex_grant4),
	.datab(!mutex_grant2),
	.datac(!master_write_data_15),
	.datad(!master_writedata_15),
	.datae(!\reg_rwdata~54_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~55 .extended_lut = "off";
defparam \reg_rwdata~55 .lut_mask = 64'hFAC80000FAC80000;
defparam \reg_rwdata~55 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~56 (
	.dataa(!sel_enabled_and_granted_0),
	.datab(!sel_enabled_and_granted_1),
	.datac(!\always2~3_combout ),
	.datad(!\l2pch|rom_l2p_ch_rtl_0|auto_generated|ram_block1a15~PORTBDATAOUT0 ),
	.datae(!reconfig_from_xcvr_15),
	.dataf(!reconfig_from_xcvr_61),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~56 .extended_lut = "off";
defparam \reg_rwdata~56 .lut_mask = 64'h000F505F303F707F;
defparam \reg_rwdata~56 .shared_arith = "off";

cyclonev_lcell_comb \reg_rwdata~57 (
	.dataa(!mutex_grant3),
	.datab(!\always2~0_combout ),
	.datac(!master_writedata_151),
	.datad(!\reg_rwdata~55_combout ),
	.datae(!\reg_rwdata~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_rwdata~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_rwdata~57 .extended_lut = "off";
defparam \reg_rwdata~57 .lut_mask = 64'h3301FFCD3301FFCD;
defparam \reg_rwdata~57 .shared_arith = "off";

cyclonev_lcell_comb \always7~0 (
	.dataa(!\always6~0_combout ),
	.datab(!wbasic_writedata_1_8),
	.datac(!wbasic_writedata_2_8),
	.datad(!wbasic_writedata_0_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always7~0 .extended_lut = "off";
defparam \always7~0 .lut_mask = 64'h4000400040004000;
defparam \always7~0 .shared_arith = "off";

cyclonev_lcell_comb \reco_write~0 (
	.dataa(!\lif_inwait~q ),
	.datab(!\reg_write_incr~q ),
	.datac(!wbasic_writedata_3_8),
	.datad(!\always2~0_combout ),
	.datae(!\always7~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_write~0 .extended_lut = "off";
defparam \reco_write~0 .lut_mask = 64'h0022F0F20022F0F2;
defparam \reco_write~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!\reg_is_phys_addr~q ),
	.datab(!\reg_addr[11]~q ),
	.datac(!\reco_addr_load_cntr[1]~q ),
	.datad(!\reco_addr_load_cntr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'h0070007000700070;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~1 (
	.dataa(!\reg_is_phys_addr~q ),
	.datab(!\reco_addr_load_cntr[1]~q ),
	.datac(!\reco_addr_load_cntr[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~1 .extended_lut = "off";
defparam \always10~1 .lut_mask = 64'h0808080808080808;
defparam \always10~1 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~2 (
	.dataa(!\reg_addr[0]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[0]~q ),
	.datae(!\Add3~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~2 .extended_lut = "off";
defparam \reco_addr~2 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~2 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~3 (
	.dataa(!\reg_addr[1]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[1]~q ),
	.datae(!\Add3~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~3 .extended_lut = "off";
defparam \reco_addr~3 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~3 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~4 (
	.dataa(!\reg_addr[2]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[2]~q ),
	.datae(!\Add3~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~4 .extended_lut = "off";
defparam \reco_addr~4 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~4 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~5 (
	.dataa(!\reg_addr[3]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[3]~q ),
	.datae(!\Add3~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~5 .extended_lut = "off";
defparam \reco_addr~5 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~5 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~6 (
	.dataa(!\reg_addr[4]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[4]~q ),
	.datae(!\Add3~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~6 .extended_lut = "off";
defparam \reco_addr~6 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~6 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~7 (
	.dataa(!\reg_addr[5]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[5]~q ),
	.datae(!\Add3~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~7 .extended_lut = "off";
defparam \reco_addr~7 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~7 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~8 (
	.dataa(!\reg_addr[6]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[6]~q ),
	.datae(!\Add3~29_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~8 .extended_lut = "off";
defparam \reco_addr~8 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~8 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~9 (
	.dataa(!\reg_addr[7]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[7]~q ),
	.datae(!\Add3~33_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~9 .extended_lut = "off";
defparam \reco_addr~9 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~9 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~10 (
	.dataa(!\reg_addr[8]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[8]~q ),
	.datae(!\Add3~37_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~10 .extended_lut = "off";
defparam \reco_addr~10 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~10 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~11 (
	.dataa(!\reg_addr[9]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[9]~q ),
	.datae(!\Add3~41_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~11 .extended_lut = "off";
defparam \reco_addr~11 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~11 .shared_arith = "off";

cyclonev_lcell_comb \reco_addr~12 (
	.dataa(!\reg_addr[10]~q ),
	.datab(!\always10~0_combout ),
	.datac(!\always10~1_combout ),
	.datad(!\l2paddr|physical_addr[10]~q ),
	.datae(!\Add3~45_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reco_addr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reco_addr~12 .extended_lut = "off";
defparam \reco_addr~12 .lut_mask = 64'h111DD1DD111DD1DD;
defparam \reco_addr~12 .shared_arith = "off";

cyclonev_lcell_comb \always6~1 (
	.dataa(!\reg_addr[0]~q ),
	.datab(!\reg_addr[1]~q ),
	.datac(!wbasic_writedata_3_8),
	.datad(!\always7~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~1 .extended_lut = "off";
defparam \always6~1 .lut_mask = 64'h0008000800080008;
defparam \always6~1 .shared_arith = "off";

cyclonev_lcell_comb \reg_plock~0 (
	.dataa(!reg_plock1),
	.datab(!wbasic_writedata_1_8),
	.datac(!wbasic_writedata_2_8),
	.datad(!wbasic_writedata_0_8),
	.datae(!wbasic_writedata_3_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_plock~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_plock~0 .extended_lut = "off";
defparam \reg_plock~0 .lut_mask = 64'h515D5555515D5555;
defparam \reg_plock~0 .shared_arith = "off";

cyclonev_lcell_comb \reg_plock~1 (
	.dataa(!reg_plock1),
	.datab(!\always2~1_combout ),
	.datac(!\lif_is_active_last~q ),
	.datad(!lif_is_active),
	.datae(!\reg_plock~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_plock~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_plock~1 .extended_lut = "off";
defparam \reg_plock~1 .lut_mask = 64'h04C437F704C437F7;
defparam \reg_plock~1 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_av_xrbasic_l2p_addr (
	ram_block1a0,
	reg_addr_0,
	reg_addr_1,
	ram_block1a1,
	reg_addr_2,
	ram_block1a2,
	reg_addr_3,
	reg_addr_4,
	reg_addr_5,
	reg_addr_6,
	reg_addr_7,
	reg_addr_8,
	reg_addr_9,
	reg_addr_10,
	reg_addr_11,
	physical_addr_11,
	physical_addr_0,
	physical_addr_1,
	physical_addr_2,
	physical_addr_3,
	physical_addr_4,
	physical_addr_5,
	physical_addr_6,
	physical_addr_7,
	physical_addr_8,
	physical_addr_9,
	physical_addr_10,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	ram_block1a0;
input 	reg_addr_0;
input 	reg_addr_1;
input 	ram_block1a1;
input 	reg_addr_2;
input 	ram_block1a2;
input 	reg_addr_3;
input 	reg_addr_4;
input 	reg_addr_5;
input 	reg_addr_6;
input 	reg_addr_7;
input 	reg_addr_8;
input 	reg_addr_9;
input 	reg_addr_10;
input 	reg_addr_11;
output 	physical_addr_11;
output 	physical_addr_0;
output 	physical_addr_1;
output 	physical_addr_2;
output 	physical_addr_3;
output 	physical_addr_4;
output 	physical_addr_5;
output 	physical_addr_6;
output 	physical_addr_7;
output 	physical_addr_8;
output 	physical_addr_9;
output 	physical_addr_10;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Decoder0~1_combout ;
wire \Decoder0~0_combout ;
wire \Add0~6 ;
wire \Add0~10 ;
wire \Add0~14 ;
wire \Add0~18 ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~30 ;
wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~9_sumout ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \Add0~29_sumout ;


dffeas \physical_addr[11] (
	.clk(mgmt_clk_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_11),
	.prn(vcc));
defparam \physical_addr[11] .is_wysiwyg = "true";
defparam \physical_addr[11] .power_up = "low";

dffeas \physical_addr[0] (
	.clk(mgmt_clk_clk),
	.d(reg_addr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_0),
	.prn(vcc));
defparam \physical_addr[0] .is_wysiwyg = "true";
defparam \physical_addr[0] .power_up = "low";

dffeas \physical_addr[1] (
	.clk(mgmt_clk_clk),
	.d(reg_addr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_1),
	.prn(vcc));
defparam \physical_addr[1] .is_wysiwyg = "true";
defparam \physical_addr[1] .power_up = "low";

dffeas \physical_addr[2] (
	.clk(mgmt_clk_clk),
	.d(reg_addr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_2),
	.prn(vcc));
defparam \physical_addr[2] .is_wysiwyg = "true";
defparam \physical_addr[2] .power_up = "low";

dffeas \physical_addr[3] (
	.clk(mgmt_clk_clk),
	.d(reg_addr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_3),
	.prn(vcc));
defparam \physical_addr[3] .is_wysiwyg = "true";
defparam \physical_addr[3] .power_up = "low";

dffeas \physical_addr[4] (
	.clk(mgmt_clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_4),
	.prn(vcc));
defparam \physical_addr[4] .is_wysiwyg = "true";
defparam \physical_addr[4] .power_up = "low";

dffeas \physical_addr[5] (
	.clk(mgmt_clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_5),
	.prn(vcc));
defparam \physical_addr[5] .is_wysiwyg = "true";
defparam \physical_addr[5] .power_up = "low";

dffeas \physical_addr[6] (
	.clk(mgmt_clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_6),
	.prn(vcc));
defparam \physical_addr[6] .is_wysiwyg = "true";
defparam \physical_addr[6] .power_up = "low";

dffeas \physical_addr[7] (
	.clk(mgmt_clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_7),
	.prn(vcc));
defparam \physical_addr[7] .is_wysiwyg = "true";
defparam \physical_addr[7] .power_up = "low";

dffeas \physical_addr[8] (
	.clk(mgmt_clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_8),
	.prn(vcc));
defparam \physical_addr[8] .is_wysiwyg = "true";
defparam \physical_addr[8] .power_up = "low";

dffeas \physical_addr[9] (
	.clk(mgmt_clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_9),
	.prn(vcc));
defparam \physical_addr[9] .is_wysiwyg = "true";
defparam \physical_addr[9] .power_up = "low";

dffeas \physical_addr[10] (
	.clk(mgmt_clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(physical_addr_10),
	.prn(vcc));
defparam \physical_addr[10] .is_wysiwyg = "true";
defparam \physical_addr[10] .power_up = "low";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!ram_block1a0),
	.datab(!ram_block1a1),
	.datac(!ram_block1a2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!ram_block1a0),
	.datab(!ram_block1a1),
	.datac(!ram_block1a2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!reg_addr_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!reg_addr_5),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reg_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!reg_addr_7),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!ram_block1a0),
	.datab(gnd),
	.datac(!ram_block1a1),
	.datad(!ram_block1a2),
	.datae(gnd),
	.dataf(!reg_addr_8),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF0000005A00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!reg_addr_9),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reg_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!reg_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~1 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_av_xrbasic_l2p_rom (
	ram_block1a0,
	ram_block1a01,
	reg_addr_0,
	reg_addr_1,
	ram_block1a1,
	ram_block1a11,
	ram_block1a2,
	ram_block1a21,
	ram_block1a3,
	ram_block1a31,
	ram_block1a16,
	ram_block1a17,
	ram_block1a18,
	ram_block1a19,
	ram_block1a20,
	ram_block1a4,
	ram_block1a211,
	ram_block1a5,
	ram_block1a22,
	ram_block1a6,
	ram_block1a23,
	ram_block1a7,
	ram_block1a24,
	ram_block1a8,
	ram_block1a25,
	ram_block1a9,
	ram_block1a26,
	ram_block1a10,
	ram_block1a27,
	ram_block1a111,
	ram_block1a28,
	ram_block1a12,
	ram_block1a29,
	ram_block1a13,
	ram_block1a30,
	ram_block1a14,
	ram_block1a311,
	ram_block1a15,
	reg_lch_0,
	reg_lch_1,
	reg_lch_2,
	reg_lch_3,
	reg_lch_4,
	GND_port,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	ram_block1a0;
output 	ram_block1a01;
input 	reg_addr_0;
input 	reg_addr_1;
output 	ram_block1a1;
output 	ram_block1a11;
output 	ram_block1a2;
output 	ram_block1a21;
output 	ram_block1a3;
output 	ram_block1a31;
output 	ram_block1a16;
output 	ram_block1a17;
output 	ram_block1a18;
output 	ram_block1a19;
output 	ram_block1a20;
output 	ram_block1a4;
output 	ram_block1a211;
output 	ram_block1a5;
output 	ram_block1a22;
output 	ram_block1a6;
output 	ram_block1a23;
output 	ram_block1a7;
output 	ram_block1a24;
output 	ram_block1a8;
output 	ram_block1a25;
output 	ram_block1a9;
output 	ram_block1a26;
output 	ram_block1a10;
output 	ram_block1a27;
output 	ram_block1a111;
output 	ram_block1a28;
output 	ram_block1a12;
output 	ram_block1a29;
output 	ram_block1a13;
output 	ram_block1a30;
output 	ram_block1a14;
output 	ram_block1a311;
output 	ram_block1a15;
input 	reg_lch_0;
input 	reg_lch_1;
input 	reg_lch_2;
input 	reg_lch_3;
input 	reg_lch_4;
input 	GND_port;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31~portadataout ;
wire \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15~portadataout ;

wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15_PORTADATAOUT_bus ;
wire [143:0] \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ;

assign ram_block1a0 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus [0];

assign ram_block1a01 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];

assign ram_block1a1 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1_PORTADATAOUT_bus [0];

assign ram_block1a11 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus [0];

assign ram_block1a2 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2_PORTADATAOUT_bus [0];

assign ram_block1a21 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus [0];

assign ram_block1a3 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3_PORTADATAOUT_bus [0];

assign ram_block1a31 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16_PORTADATAOUT_bus [0];

assign ram_block1a16 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17_PORTADATAOUT_bus [0];

assign ram_block1a17 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18_PORTADATAOUT_bus [0];

assign ram_block1a18 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19_PORTADATAOUT_bus [0];

assign ram_block1a19 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20_PORTADATAOUT_bus [0];

assign ram_block1a20 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus [0];

assign ram_block1a4 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21_PORTADATAOUT_bus [0];

assign ram_block1a211 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5_PORTADATAOUT_bus [0];

assign ram_block1a5 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22_PORTADATAOUT_bus [0];

assign ram_block1a22 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6_PORTADATAOUT_bus [0];

assign ram_block1a6 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23_PORTADATAOUT_bus [0];

assign ram_block1a23 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7_PORTADATAOUT_bus [0];

assign ram_block1a7 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24_PORTADATAOUT_bus [0];

assign ram_block1a24 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8_PORTADATAOUT_bus [0];

assign ram_block1a8 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25_PORTADATAOUT_bus [0];

assign ram_block1a25 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9_PORTADATAOUT_bus [0];

assign ram_block1a9 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26_PORTADATAOUT_bus [0];

assign ram_block1a26 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10_PORTADATAOUT_bus [0];

assign ram_block1a10 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27_PORTADATAOUT_bus [0];

assign ram_block1a27 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11_PORTADATAOUT_bus [0];

assign ram_block1a111 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28_PORTADATAOUT_bus [0];

assign ram_block1a28 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus [0];

assign ram_block1a12 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29_PORTADATAOUT_bus [0];

assign ram_block1a29 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13_PORTADATAOUT_bus [0];

assign ram_block1a13 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30_PORTADATAOUT_bus [0];

assign ram_block1a30 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14_PORTADATAOUT_bus [0];

assign ram_block1a14 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31_PORTADATAOUT_bus [0];

assign ram_block1a311 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus [0];

assign \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15~portadataout  = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15_PORTADATAOUT_bus [0];

assign ram_block1a15 = \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus [0];

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_first_bit_number = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a0 .mem_init0 = "11111111111111111111111111111100";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a1_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_first_bit_number = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_first_bit_number = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a1 .mem_init0 = "11111111111111111111111111111100";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a2_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_first_bit_number = 2;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_first_bit_number = 2;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a2 .mem_init0 = "11111111111111111111111111111100";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a3_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_first_bit_number = 3;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_first_bit_number = 3;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a3 .mem_init0 = "11111111111111111111111111111110";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a16_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_first_bit_number = 16;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_first_bit_number = 16;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a16 .mem_init0 = "22222222222222222222222222222222";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a17_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_first_bit_number = 17;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_first_bit_number = 17;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a17 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a18_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_first_bit_number = 18;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_first_bit_number = 18;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a18 .mem_init0 = "44444444444444444444444444444444";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a19_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_first_bit_number = 19;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_first_bit_number = 19;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a19 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a20_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_first_bit_number = 20;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_first_bit_number = 20;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a20 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_first_bit_number = 4;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a4 .mem_init0 = "44444444444444444444444444444444";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a21_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_first_bit_number = 21;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_first_bit_number = 21;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a21 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a5_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_first_bit_number = 5;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_first_bit_number = 5;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a5 .mem_init0 = "22222222222222222222222222222222";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a22_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_first_bit_number = 22;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_first_bit_number = 22;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a22 .mem_init0 = "22222222222222222222222222222222";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a6_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_first_bit_number = 6;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_first_bit_number = 6;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a6 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a23_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_first_bit_number = 23;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_first_bit_number = 23;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a23 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a7_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_first_bit_number = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_first_bit_number = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a7 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a24_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_first_bit_number = 24;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_first_bit_number = 24;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a24 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a8_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_first_bit_number = 8;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_first_bit_number = 8;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a8 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a25_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_first_bit_number = 25;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_first_bit_number = 25;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a25 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a9_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_first_bit_number = 9;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_first_bit_number = 9;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a9 .mem_init0 = "44444444444444444444444444444444";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a26_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_first_bit_number = 26;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_first_bit_number = 26;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a26 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a10_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_first_bit_number = 10;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_first_bit_number = 10;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a10 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a27_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_first_bit_number = 27;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_first_bit_number = 27;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a27 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a11_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_first_bit_number = 11;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_first_bit_number = 11;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a11 .mem_init0 = "22222222222222222222222222222222";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a28_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_first_bit_number = 28;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_first_bit_number = 28;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a28 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_first_bit_number = 12;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_first_bit_number = 12;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a12 .mem_init0 = "44444444444444444444444444444444";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a29_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_first_bit_number = 29;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_first_bit_number = 29;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a29 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a13_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_first_bit_number = 13;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_first_bit_number = 13;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a13 .mem_init0 = "44444444444444444444444444444444";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a30_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_first_bit_number = 30;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_first_bit_number = 30;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a30 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a14_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_first_bit_number = 14;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_first_bit_number = 14;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a14 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a31_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_first_bit_number = 31;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_first_bit_number = 31;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a31 .mem_init0 = "00000000000000000000000000000000";

cyclonev_ram_block \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 (
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mgmt_clk_clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,GND_port,GND_port}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,reg_lch_4,reg_lch_3,reg_lch_2,reg_lch_1,reg_lch_0,reg_addr_1,reg_addr_0}),
	.portbbyteenamasks(1'b1),
	.portadataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a15_PORTADATAOUT_bus ),
	.portbdataout(\rom_l2p_ch_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .data_interleave_offset_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .data_interleave_width_in_bits = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .init_file = "db/RECONFIGURE_IP.ram0_av_xrbasic_l2p_rom_f62b5f4.hdl.mif";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .init_file_layout = "port_a";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .logical_ram_name = "alt_xcvr_reconfig:reconfigure_ip_inst|alt_xcvr_reconfig_basic:basic|av_xcvr_reconfig_basic:a5|av_xrbasic_lif:lif[0].logical_if|av_xrbasic_lif_csr:lif_csr|av_xrbasic_l2p_rom:l2pch|altsyncram:rom_l2p_ch_rtl_0|altsyncram_0l22:auto_generated|ALTSYNCRAM";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .mixed_port_feed_through_mode = "dont_care";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .operation_mode = "bidir_dual_port";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_first_bit_number = 15;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_address_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_address_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_address_width = 7;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_data_in_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clear = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clock = "none";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_data_width = 1;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_first_address = 0;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_first_bit_number = 15;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_last_address = 127;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_depth = 128;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_width = 32;
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_read_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .port_b_write_enable_clock = "clock0";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .ram_block_type = "M20K";
defparam \rom_l2p_ch_rtl_0|auto_generated|ram_block1a15 .mem_init0 = "22222222222222222222222222222222";

endmodule

module RECONFIGURE_IP_csr_mux (
	ram_block1a0,
	ram_block1a1,
	ram_block1a2,
	pif_enabled_and_granted_0,
	pif_enabled_and_granted_1,
	pif_testbus_groups_0_1,
	pif_testbus_groups_16_1,
	out_narrow_0,
	pif_testbus_groups_1_1,
	pif_testbus_groups_17_1,
	out_narrow_1,
	pif_testbus_groups_2_1,
	pif_testbus_groups_18_1,
	out_narrow_2,
	pif_testbus_groups_3_1,
	pif_testbus_groups_19_1,
	out_narrow_3,
	reconfig_from_xcvr_24,
	reconfig_from_xcvr_70,
	reconfig_from_xcvr_25,
	reconfig_from_xcvr_71,
	reconfig_from_xcvr_26,
	reconfig_from_xcvr_72,
	reconfig_from_xcvr_27,
	reconfig_from_xcvr_73)/* synthesis synthesis_greybox=0 */;
input 	ram_block1a0;
input 	ram_block1a1;
input 	ram_block1a2;
input 	pif_enabled_and_granted_0;
input 	pif_enabled_and_granted_1;
input 	pif_testbus_groups_0_1;
input 	pif_testbus_groups_16_1;
output 	out_narrow_0;
input 	pif_testbus_groups_1_1;
input 	pif_testbus_groups_17_1;
output 	out_narrow_1;
input 	pif_testbus_groups_2_1;
input 	pif_testbus_groups_18_1;
output 	out_narrow_2;
input 	pif_testbus_groups_3_1;
input 	pif_testbus_groups_19_1;
output 	out_narrow_3;
input 	reconfig_from_xcvr_24;
input 	reconfig_from_xcvr_70;
input 	reconfig_from_xcvr_25;
input 	reconfig_from_xcvr_71;
input 	reconfig_from_xcvr_26;
input 	reconfig_from_xcvr_72;
input 	reconfig_from_xcvr_27;
input 	reconfig_from_xcvr_73;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_narrow[0]~8_combout ;
wire \out_narrow[0]~1_combout ;
wire \out_narrow[0]~0_combout ;
wire \out_narrow[1]~10_combout ;
wire \out_narrow[1]~3_combout ;
wire \out_narrow[1]~2_combout ;
wire \out_narrow[2]~12_combout ;
wire \out_narrow[2]~5_combout ;
wire \out_narrow[2]~4_combout ;
wire \out_narrow[3]~14_combout ;
wire \out_narrow[3]~7_combout ;
wire \out_narrow[3]~6_combout ;


cyclonev_lcell_comb \out_narrow[0] (
	.dataa(!ram_block1a2),
	.datab(!\out_narrow[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_narrow_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[0] .extended_lut = "off";
defparam \out_narrow[0] .lut_mask = 64'h2222222222222222;
defparam \out_narrow[0] .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[1] (
	.dataa(!ram_block1a2),
	.datab(!\out_narrow[1]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_narrow_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[1] .extended_lut = "off";
defparam \out_narrow[1] .lut_mask = 64'h2222222222222222;
defparam \out_narrow[1] .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[2] (
	.dataa(!ram_block1a2),
	.datab(!\out_narrow[2]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_narrow_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[2] .extended_lut = "off";
defparam \out_narrow[2] .lut_mask = 64'h2222222222222222;
defparam \out_narrow[2] .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[3] (
	.dataa(!ram_block1a2),
	.datab(!\out_narrow[3]~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_narrow_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[3] .extended_lut = "off";
defparam \out_narrow[3] .lut_mask = 64'h2222222222222222;
defparam \out_narrow[3] .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[0]~8 (
	.dataa(!pif_enabled_and_granted_0),
	.datab(!pif_enabled_and_granted_1),
	.datac(!ram_block1a1),
	.datad(!reconfig_from_xcvr_24),
	.datae(!reconfig_from_xcvr_70),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[0]~8 .extended_lut = "off";
defparam \out_narrow[0]~8 .lut_mask = 64'h0050307000503070;
defparam \out_narrow[0]~8 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[0]~1 (
	.dataa(!pif_testbus_groups_0_1),
	.datab(!pif_testbus_groups_16_1),
	.datac(!ram_block1a1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[0]~1 .extended_lut = "off";
defparam \out_narrow[0]~1 .lut_mask = 64'hACACACACACACACAC;
defparam \out_narrow[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[0]~0 (
	.dataa(!\out_narrow[0]~8_combout ),
	.datab(!\out_narrow[0]~1_combout ),
	.datac(!ram_block1a0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[0]~0 .extended_lut = "off";
defparam \out_narrow[0]~0 .lut_mask = 64'hC5C5C5C5C5C5C5C5;
defparam \out_narrow[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[1]~10 (
	.dataa(!pif_enabled_and_granted_0),
	.datab(!pif_enabled_and_granted_1),
	.datac(!ram_block1a1),
	.datad(!reconfig_from_xcvr_25),
	.datae(!reconfig_from_xcvr_71),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[1]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[1]~10 .extended_lut = "off";
defparam \out_narrow[1]~10 .lut_mask = 64'h0050307000503070;
defparam \out_narrow[1]~10 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[1]~3 (
	.dataa(!pif_testbus_groups_1_1),
	.datab(!pif_testbus_groups_17_1),
	.datac(!ram_block1a1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[1]~3 .extended_lut = "off";
defparam \out_narrow[1]~3 .lut_mask = 64'hACACACACACACACAC;
defparam \out_narrow[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[1]~2 (
	.dataa(!\out_narrow[1]~10_combout ),
	.datab(!\out_narrow[1]~3_combout ),
	.datac(!ram_block1a0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[1]~2 .extended_lut = "off";
defparam \out_narrow[1]~2 .lut_mask = 64'hC5C5C5C5C5C5C5C5;
defparam \out_narrow[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[2]~12 (
	.dataa(!pif_enabled_and_granted_0),
	.datab(!pif_enabled_and_granted_1),
	.datac(!ram_block1a1),
	.datad(!reconfig_from_xcvr_26),
	.datae(!reconfig_from_xcvr_72),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[2]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[2]~12 .extended_lut = "off";
defparam \out_narrow[2]~12 .lut_mask = 64'h0050307000503070;
defparam \out_narrow[2]~12 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[2]~5 (
	.dataa(!pif_testbus_groups_2_1),
	.datab(!pif_testbus_groups_18_1),
	.datac(!ram_block1a1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[2]~5 .extended_lut = "off";
defparam \out_narrow[2]~5 .lut_mask = 64'hACACACACACACACAC;
defparam \out_narrow[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[2]~4 (
	.dataa(!\out_narrow[2]~12_combout ),
	.datab(!\out_narrow[2]~5_combout ),
	.datac(!ram_block1a0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[2]~4 .extended_lut = "off";
defparam \out_narrow[2]~4 .lut_mask = 64'hC5C5C5C5C5C5C5C5;
defparam \out_narrow[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[3]~14 (
	.dataa(!pif_enabled_and_granted_0),
	.datab(!pif_enabled_and_granted_1),
	.datac(!ram_block1a1),
	.datad(!reconfig_from_xcvr_27),
	.datae(!reconfig_from_xcvr_73),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[3]~14 .extended_lut = "off";
defparam \out_narrow[3]~14 .lut_mask = 64'h0050307000503070;
defparam \out_narrow[3]~14 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[3]~7 (
	.dataa(!pif_testbus_groups_3_1),
	.datab(!pif_testbus_groups_19_1),
	.datac(!ram_block1a1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[3]~7 .extended_lut = "off";
defparam \out_narrow[3]~7 .lut_mask = 64'hACACACACACACACAC;
defparam \out_narrow[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \out_narrow[3]~6 (
	.dataa(!\out_narrow[3]~14_combout ),
	.datab(!\out_narrow[3]~7_combout ),
	.datac(!ram_block1a0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_narrow[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_narrow[3]~6 .extended_lut = "off";
defparam \out_narrow[3]~6 .lut_mask = 64'hC5C5C5C5C5C5C5C5;
defparam \out_narrow[3]~6 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_cal_seq (
	reconfig_busy1,
	offset_cancellation_done,
	tx_cal_busy1,
	rx_cal_busy1,
	uif_busy,
	pll_mif_busy,
	stateSTATE_IDLE,
	ifsel_notdone_resync,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	reconfig_busy1;
input 	offset_cancellation_done;
output 	tx_cal_busy1;
output 	rx_cal_busy1;
input 	uif_busy;
input 	pll_mif_busy;
input 	stateSTATE_IDLE;
input 	ifsel_notdone_resync;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~combout ;
wire \rx_cal_busy~0_combout ;


dffeas reconfig_busy(
	.clk(mgmt_clk_clk),
	.d(\WideOr0~combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reconfig_busy1),
	.prn(vcc));
defparam reconfig_busy.is_wysiwyg = "true";
defparam reconfig_busy.power_up = "low";

dffeas tx_cal_busy(
	.clk(mgmt_clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_cal_busy1),
	.prn(vcc));
defparam tx_cal_busy.is_wysiwyg = "true";
defparam tx_cal_busy.power_up = "low";

dffeas rx_cal_busy(
	.clk(mgmt_clk_clk),
	.d(\rx_cal_busy~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rx_cal_busy1),
	.prn(vcc));
defparam rx_cal_busy.is_wysiwyg = "true";
defparam rx_cal_busy.power_up = "low";

cyclonev_lcell_comb WideOr0(
	.dataa(!offset_cancellation_done),
	.datab(!uif_busy),
	.datac(!pll_mif_busy),
	.datad(!stateSTATE_IDLE),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h4000400040004000;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \rx_cal_busy~0 (
	.dataa(!offset_cancellation_done),
	.datab(!rx_cal_busy1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_cal_busy~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_cal_busy~0 .extended_lut = "off";
defparam \rx_cal_busy~0 .lut_mask = 64'h7777777777777777;
defparam \rx_cal_busy~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_direct (
	Equal2,
	reg_arb_req1,
	grant_4,
	mutex_grant,
	basic_write,
	reset,
	master_read,
	reconfig_mgmt_address_3,
	reconfig_mgmt_address_4,
	reconfig_mgmt_address_5,
	reconfig_mgmt_address_6,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	clk,
	reconfig_mgmt_writedata_0)/* synthesis synthesis_greybox=0 */;
input 	Equal2;
output 	reg_arb_req1;
input 	grant_4;
output 	mutex_grant;
output 	basic_write;
input 	reset;
output 	master_read;
input 	reconfig_mgmt_address_3;
input 	reconfig_mgmt_address_4;
input 	reconfig_mgmt_address_5;
input 	reconfig_mgmt_address_6;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	clk;
input 	reconfig_mgmt_writedata_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \reg_arb_req~0_combout ;


RECONFIGURE_IP_alt_arbiter_acq_1 mutex_inst(
	.reg_arb_req(reg_arb_req1),
	.grant_4(grant_4),
	.mutex_grant1(mutex_grant),
	.master_write(basic_write),
	.master_read1(master_read),
	.reconfig_mgmt_address_3(reconfig_mgmt_address_3),
	.reconfig_mgmt_address_4(reconfig_mgmt_address_4),
	.reconfig_mgmt_address_5(reconfig_mgmt_address_5),
	.reconfig_mgmt_address_6(reconfig_mgmt_address_6),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read));

dffeas reg_arb_req(
	.clk(clk),
	.d(\reg_arb_req~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reg_arb_req1),
	.prn(vcc));
defparam reg_arb_req.is_wysiwyg = "true";
defparam reg_arb_req.power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!reconfig_mgmt_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0080008000800080;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \reg_arb_req~0 (
	.dataa(!Equal2),
	.datab(!reg_arb_req1),
	.datac(!reconfig_mgmt_writedata_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reg_arb_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_arb_req~0 .extended_lut = "off";
defparam \reg_arb_req~0 .lut_mask = 64'h3327332733273327;
defparam \reg_arb_req~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_arbiter_acq_1 (
	reg_arb_req,
	grant_4,
	mutex_grant1,
	master_write,
	master_read1,
	reconfig_mgmt_address_3,
	reconfig_mgmt_address_4,
	reconfig_mgmt_address_5,
	reconfig_mgmt_address_6,
	reconfig_mgmt_write,
	reconfig_mgmt_read)/* synthesis synthesis_greybox=0 */;
input 	reg_arb_req;
input 	grant_4;
output 	mutex_grant1;
output 	master_write;
output 	master_read1;
input 	reconfig_mgmt_address_3;
input 	reconfig_mgmt_address_4;
input 	reconfig_mgmt_address_5;
input 	reconfig_mgmt_address_6;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb mutex_grant(
	.dataa(!reg_arb_req),
	.datab(!grant_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mutex_grant1),
	.sumout(),
	.cout(),
	.shareout());
defparam mutex_grant.extended_lut = "off";
defparam mutex_grant.lut_mask = 64'h1111111111111111;
defparam mutex_grant.shared_arith = "off";

cyclonev_lcell_comb \master_write~0 (
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!mutex_grant1),
	.dataf(!reconfig_mgmt_write),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write~0 .extended_lut = "off";
defparam \master_write~0 .lut_mask = 64'h0000000000000800;
defparam \master_write~0 .shared_arith = "off";

cyclonev_lcell_comb master_read(
	.dataa(!reconfig_mgmt_address_3),
	.datab(!reconfig_mgmt_address_4),
	.datac(!reconfig_mgmt_address_5),
	.datad(!reconfig_mgmt_address_6),
	.datae(!reconfig_mgmt_read),
	.dataf(!mutex_grant1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_read1),
	.sumout(),
	.cout(),
	.shareout());
defparam master_read.extended_lut = "off";
defparam master_read.lut_mask = 64'h0000000000000800;
defparam master_read.shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_mif (
	user_reconfig_readdata_12,
	basic_reconfig_readdata_12,
	user_reconfig_readdata_13,
	basic_reconfig_readdata_13,
	user_reconfig_readdata_14,
	basic_reconfig_readdata_14,
	user_reconfig_readdata_15,
	basic_reconfig_readdata_15,
	user_reconfig_readdata_16,
	basic_reconfig_readdata_16,
	user_reconfig_readdata_17,
	basic_reconfig_readdata_17,
	user_reconfig_readdata_18,
	basic_reconfig_readdata_18,
	user_reconfig_readdata_19,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	user_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	user_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	user_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	user_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	user_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	user_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	user_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	user_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	user_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	user_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	user_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	user_reconfig_readdata_31,
	stream_address_0,
	stream_address_1,
	stream_address_2,
	stream_address_3,
	stream_address_4,
	stream_address_5,
	stream_address_6,
	stream_address_7,
	stream_address_8,
	stream_address_9,
	stream_address_10,
	stream_address_11,
	stream_address_12,
	stream_address_13,
	stream_address_14,
	stream_address_15,
	stream_address_16,
	stream_address_17,
	stream_address_18,
	stream_address_19,
	stream_address_20,
	stream_address_21,
	stream_address_22,
	stream_address_23,
	stream_address_24,
	stream_address_25,
	stream_address_26,
	stream_address_27,
	stream_address_28,
	stream_address_29,
	stream_address_30,
	stream_address_31,
	user_reconfig_readdata_0,
	Equal3,
	basic_reconfig_readdata_0,
	user_reconfig_readdata_1,
	basic_reconfig_readdata_1,
	user_reconfig_readdata_2,
	basic_reconfig_readdata_2,
	user_reconfig_readdata_3,
	basic_reconfig_readdata_3,
	user_reconfig_readdata_4,
	basic_reconfig_readdata_4,
	user_reconfig_readdata_5,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	user_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	user_reconfig_readdata_7,
	reconfig_mgmt_readdata_8,
	basic_reconfig_readdata_8,
	user_reconfig_readdata_8,
	user_reconfig_readdata_9,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	user_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	user_reconfig_readdata_11,
	master_write,
	grant_7,
	mutex_req,
	mutex_grant,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	stream_read,
	uif_busy,
	pll_mif_busy,
	ifsel_notdone_resync,
	uif_logical_ch_addr_0,
	comb,
	uif_logical_ch_addr_1,
	uif_logical_ch_addr_2,
	uif_logical_ch_addr_3,
	user_reconfig_readdata_101,
	uif_logical_ch_addr_4,
	uif_logical_ch_addr_5,
	uif_logical_ch_addr_6,
	uif_logical_ch_addr_7,
	uif_logical_ch_addr_8,
	uif_logical_ch_addr_9,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	pll_go,
	uif_mode_0,
	Mux0,
	Mux3,
	WideOr0,
	pll_type,
	mif_rec_addr_7,
	mif_rec_addr_5,
	mif_rec_addr_6,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mif_waitrequest,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15,
	reconfig_mif_readdata_15,
	reconfig_mif_readdata_14,
	reconfig_mif_readdata_13,
	reconfig_mif_readdata_12,
	reconfig_mif_readdata_11,
	reconfig_mif_readdata_1,
	reconfig_mif_readdata_0,
	reconfig_mif_readdata_4,
	reconfig_mif_readdata_3,
	reconfig_mif_readdata_2,
	reconfig_mif_readdata_7,
	reconfig_mif_readdata_5,
	reconfig_mif_readdata_6,
	reconfig_mif_readdata_8,
	reconfig_mif_readdata_9,
	reconfig_mif_readdata_10)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_12;
input 	basic_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
input 	basic_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
input 	basic_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
input 	basic_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
input 	basic_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
input 	basic_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
input 	basic_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
output 	user_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
output 	user_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
output 	user_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
output 	user_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
output 	user_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
output 	user_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
output 	user_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
output 	user_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
output 	user_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
output 	user_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
output 	user_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	user_reconfig_readdata_31;
output 	stream_address_0;
output 	stream_address_1;
output 	stream_address_2;
output 	stream_address_3;
output 	stream_address_4;
output 	stream_address_5;
output 	stream_address_6;
output 	stream_address_7;
output 	stream_address_8;
output 	stream_address_9;
output 	stream_address_10;
output 	stream_address_11;
output 	stream_address_12;
output 	stream_address_13;
output 	stream_address_14;
output 	stream_address_15;
output 	stream_address_16;
output 	stream_address_17;
output 	stream_address_18;
output 	stream_address_19;
output 	stream_address_20;
output 	stream_address_21;
output 	stream_address_22;
output 	stream_address_23;
output 	stream_address_24;
output 	stream_address_25;
output 	stream_address_26;
output 	stream_address_27;
output 	stream_address_28;
output 	stream_address_29;
output 	stream_address_30;
output 	stream_address_31;
output 	user_reconfig_readdata_0;
input 	Equal3;
input 	basic_reconfig_readdata_0;
output 	user_reconfig_readdata_1;
input 	basic_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
input 	basic_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
input 	basic_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
input 	basic_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
output 	user_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
output 	user_reconfig_readdata_7;
input 	reconfig_mgmt_readdata_8;
input 	basic_reconfig_readdata_8;
output 	user_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
output 	user_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	user_reconfig_readdata_11;
output 	master_write;
input 	grant_7;
output 	mutex_req;
output 	mutex_grant;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
output 	stream_read;
output 	uif_busy;
input 	pll_mif_busy;
input 	ifsel_notdone_resync;
output 	uif_logical_ch_addr_0;
input 	comb;
output 	uif_logical_ch_addr_1;
output 	uif_logical_ch_addr_2;
output 	uif_logical_ch_addr_3;
input 	user_reconfig_readdata_101;
output 	uif_logical_ch_addr_4;
output 	uif_logical_ch_addr_5;
output 	uif_logical_ch_addr_6;
output 	uif_logical_ch_addr_7;
output 	uif_logical_ch_addr_8;
output 	uif_logical_ch_addr_9;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
output 	pll_go;
input 	uif_mode_0;
input 	Mux0;
input 	Mux3;
input 	WideOr0;
output 	pll_type;
output 	mif_rec_addr_7;
output 	mif_rec_addr_5;
output 	mif_rec_addr_6;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mif_waitrequest;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;
input 	reconfig_mif_readdata_15;
input 	reconfig_mif_readdata_14;
input 	reconfig_mif_readdata_13;
input 	reconfig_mif_readdata_12;
input 	reconfig_mif_readdata_11;
input 	reconfig_mif_readdata_1;
input 	reconfig_mif_readdata_0;
input 	reconfig_mif_readdata_4;
input 	reconfig_mif_readdata_3;
input 	reconfig_mif_readdata_2;
input 	reconfig_mif_readdata_7;
input 	reconfig_mif_readdata_5;
input 	reconfig_mif_readdata_6;
input 	reconfig_mif_readdata_8;
input 	reconfig_mif_readdata_9;
input 	reconfig_mif_readdata_10;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



RECONFIGURE_IP_av_xcvr_reconfig_mif mif_strm_av(
	.user_reconfig_readdata_12(user_reconfig_readdata_12),
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.user_reconfig_readdata_13(user_reconfig_readdata_13),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.user_reconfig_readdata_14(user_reconfig_readdata_14),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.user_reconfig_readdata_15(user_reconfig_readdata_15),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.user_reconfig_readdata_16(user_reconfig_readdata_16),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.user_reconfig_readdata_17(user_reconfig_readdata_17),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.user_reconfig_readdata_18(user_reconfig_readdata_18),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.user_reconfig_readdata_19(user_reconfig_readdata_19),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.user_reconfig_readdata_20(user_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.user_reconfig_readdata_21(user_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.user_reconfig_readdata_22(user_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.user_reconfig_readdata_23(user_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.user_reconfig_readdata_24(user_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.user_reconfig_readdata_25(user_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.user_reconfig_readdata_26(user_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.user_reconfig_readdata_27(user_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.user_reconfig_readdata_28(user_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.user_reconfig_readdata_29(user_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.user_reconfig_readdata_30(user_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.user_reconfig_readdata_31(user_reconfig_readdata_31),
	.stream_address_0(stream_address_0),
	.stream_address_1(stream_address_1),
	.stream_address_2(stream_address_2),
	.stream_address_3(stream_address_3),
	.stream_address_4(stream_address_4),
	.stream_address_5(stream_address_5),
	.stream_address_6(stream_address_6),
	.stream_address_7(stream_address_7),
	.stream_address_8(stream_address_8),
	.stream_address_9(stream_address_9),
	.stream_address_10(stream_address_10),
	.stream_address_11(stream_address_11),
	.stream_address_12(stream_address_12),
	.stream_address_13(stream_address_13),
	.stream_address_14(stream_address_14),
	.stream_address_15(stream_address_15),
	.stream_address_16(stream_address_16),
	.stream_address_17(stream_address_17),
	.stream_address_18(stream_address_18),
	.stream_address_19(stream_address_19),
	.stream_address_20(stream_address_20),
	.stream_address_21(stream_address_21),
	.stream_address_22(stream_address_22),
	.stream_address_23(stream_address_23),
	.stream_address_24(stream_address_24),
	.stream_address_25(stream_address_25),
	.stream_address_26(stream_address_26),
	.stream_address_27(stream_address_27),
	.stream_address_28(stream_address_28),
	.stream_address_29(stream_address_29),
	.stream_address_30(stream_address_30),
	.stream_address_31(stream_address_31),
	.user_reconfig_readdata_0(user_reconfig_readdata_0),
	.Equal3(Equal3),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.user_reconfig_readdata_1(user_reconfig_readdata_1),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.user_reconfig_readdata_2(user_reconfig_readdata_2),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.user_reconfig_readdata_3(user_reconfig_readdata_3),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.user_reconfig_readdata_4(user_reconfig_readdata_4),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.user_reconfig_readdata_5(user_reconfig_readdata_5),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.user_reconfig_readdata_6(user_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.user_reconfig_readdata_7(user_reconfig_readdata_7),
	.reconfig_mgmt_readdata_8(reconfig_mgmt_readdata_8),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.user_reconfig_readdata_8(user_reconfig_readdata_8),
	.user_reconfig_readdata_9(user_reconfig_readdata_9),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.user_reconfig_readdata_10(user_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.user_reconfig_readdata_11(user_reconfig_readdata_11),
	.master_write(master_write),
	.grant_7(grant_7),
	.mutex_req(mutex_req),
	.mutex_grant(mutex_grant),
	.master_address_2(master_address_2),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg(launch_reg),
	.wait_reg(wait_reg),
	.stream_read(stream_read),
	.uif_busy(uif_busy),
	.pll_mif_busy(pll_mif_busy),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.uif_logical_ch_addr_0(uif_logical_ch_addr_0),
	.comb(comb),
	.uif_logical_ch_addr_1(uif_logical_ch_addr_1),
	.uif_logical_ch_addr_2(uif_logical_ch_addr_2),
	.uif_logical_ch_addr_3(uif_logical_ch_addr_3),
	.user_reconfig_readdata_101(user_reconfig_readdata_101),
	.uif_logical_ch_addr_4(uif_logical_ch_addr_4),
	.uif_logical_ch_addr_5(uif_logical_ch_addr_5),
	.uif_logical_ch_addr_6(uif_logical_ch_addr_6),
	.uif_logical_ch_addr_7(uif_logical_ch_addr_7),
	.uif_logical_ch_addr_8(uif_logical_ch_addr_8),
	.uif_logical_ch_addr_9(uif_logical_ch_addr_9),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.master_writedata_11(master_writedata_11),
	.master_writedata_12(master_writedata_12),
	.master_writedata_13(master_writedata_13),
	.master_writedata_14(master_writedata_14),
	.master_writedata_15(master_writedata_15),
	.pll_go(pll_go),
	.uif_mode_0(uif_mode_0),
	.Mux0(Mux0),
	.Mux3(Mux3),
	.WideOr0(WideOr0),
	.pll_type(pll_type),
	.mif_rec_addr_7(mif_rec_addr_7),
	.mif_rec_addr_5(mif_rec_addr_5),
	.mif_rec_addr_6(mif_rec_addr_6),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mif_waitrequest(reconfig_mif_waitrequest),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15),
	.reconfig_mif_readdata_15(reconfig_mif_readdata_15),
	.reconfig_mif_readdata_14(reconfig_mif_readdata_14),
	.reconfig_mif_readdata_13(reconfig_mif_readdata_13),
	.reconfig_mif_readdata_12(reconfig_mif_readdata_12),
	.reconfig_mif_readdata_11(reconfig_mif_readdata_11),
	.reconfig_mif_readdata_1(reconfig_mif_readdata_1),
	.reconfig_mif_readdata_0(reconfig_mif_readdata_0),
	.reconfig_mif_readdata_4(reconfig_mif_readdata_4),
	.reconfig_mif_readdata_3(reconfig_mif_readdata_3),
	.reconfig_mif_readdata_2(reconfig_mif_readdata_2),
	.reconfig_mif_readdata_7(reconfig_mif_readdata_7),
	.reconfig_mif_readdata_5(reconfig_mif_readdata_5),
	.reconfig_mif_readdata_6(reconfig_mif_readdata_6),
	.reconfig_mif_readdata_8(reconfig_mif_readdata_8),
	.reconfig_mif_readdata_9(reconfig_mif_readdata_9),
	.reconfig_mif_readdata_10(reconfig_mif_readdata_10));

endmodule

module RECONFIGURE_IP_av_xcvr_reconfig_mif (
	user_reconfig_readdata_12,
	basic_reconfig_readdata_12,
	user_reconfig_readdata_13,
	basic_reconfig_readdata_13,
	user_reconfig_readdata_14,
	basic_reconfig_readdata_14,
	user_reconfig_readdata_15,
	basic_reconfig_readdata_15,
	user_reconfig_readdata_16,
	basic_reconfig_readdata_16,
	user_reconfig_readdata_17,
	basic_reconfig_readdata_17,
	user_reconfig_readdata_18,
	basic_reconfig_readdata_18,
	user_reconfig_readdata_19,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	user_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	user_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	user_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	user_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	user_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	user_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	user_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	user_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	user_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	user_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	user_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	user_reconfig_readdata_31,
	stream_address_0,
	stream_address_1,
	stream_address_2,
	stream_address_3,
	stream_address_4,
	stream_address_5,
	stream_address_6,
	stream_address_7,
	stream_address_8,
	stream_address_9,
	stream_address_10,
	stream_address_11,
	stream_address_12,
	stream_address_13,
	stream_address_14,
	stream_address_15,
	stream_address_16,
	stream_address_17,
	stream_address_18,
	stream_address_19,
	stream_address_20,
	stream_address_21,
	stream_address_22,
	stream_address_23,
	stream_address_24,
	stream_address_25,
	stream_address_26,
	stream_address_27,
	stream_address_28,
	stream_address_29,
	stream_address_30,
	stream_address_31,
	user_reconfig_readdata_0,
	Equal3,
	basic_reconfig_readdata_0,
	user_reconfig_readdata_1,
	basic_reconfig_readdata_1,
	user_reconfig_readdata_2,
	basic_reconfig_readdata_2,
	user_reconfig_readdata_3,
	basic_reconfig_readdata_3,
	user_reconfig_readdata_4,
	basic_reconfig_readdata_4,
	user_reconfig_readdata_5,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	user_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	user_reconfig_readdata_7,
	reconfig_mgmt_readdata_8,
	basic_reconfig_readdata_8,
	user_reconfig_readdata_8,
	user_reconfig_readdata_9,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	user_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	user_reconfig_readdata_11,
	master_write,
	grant_7,
	mutex_req,
	mutex_grant,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	stream_read,
	uif_busy,
	pll_mif_busy,
	ifsel_notdone_resync,
	uif_logical_ch_addr_0,
	comb,
	uif_logical_ch_addr_1,
	uif_logical_ch_addr_2,
	uif_logical_ch_addr_3,
	user_reconfig_readdata_101,
	uif_logical_ch_addr_4,
	uif_logical_ch_addr_5,
	uif_logical_ch_addr_6,
	uif_logical_ch_addr_7,
	uif_logical_ch_addr_8,
	uif_logical_ch_addr_9,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	pll_go,
	uif_mode_0,
	Mux0,
	Mux3,
	WideOr0,
	pll_type,
	mif_rec_addr_7,
	mif_rec_addr_5,
	mif_rec_addr_6,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mif_waitrequest,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15,
	reconfig_mif_readdata_15,
	reconfig_mif_readdata_14,
	reconfig_mif_readdata_13,
	reconfig_mif_readdata_12,
	reconfig_mif_readdata_11,
	reconfig_mif_readdata_1,
	reconfig_mif_readdata_0,
	reconfig_mif_readdata_4,
	reconfig_mif_readdata_3,
	reconfig_mif_readdata_2,
	reconfig_mif_readdata_7,
	reconfig_mif_readdata_5,
	reconfig_mif_readdata_6,
	reconfig_mif_readdata_8,
	reconfig_mif_readdata_9,
	reconfig_mif_readdata_10)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_12;
input 	basic_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
input 	basic_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
input 	basic_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
input 	basic_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
input 	basic_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
input 	basic_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
input 	basic_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
output 	user_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
output 	user_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
output 	user_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
output 	user_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
output 	user_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
output 	user_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
output 	user_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
output 	user_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
output 	user_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
output 	user_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
output 	user_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	user_reconfig_readdata_31;
output 	stream_address_0;
output 	stream_address_1;
output 	stream_address_2;
output 	stream_address_3;
output 	stream_address_4;
output 	stream_address_5;
output 	stream_address_6;
output 	stream_address_7;
output 	stream_address_8;
output 	stream_address_9;
output 	stream_address_10;
output 	stream_address_11;
output 	stream_address_12;
output 	stream_address_13;
output 	stream_address_14;
output 	stream_address_15;
output 	stream_address_16;
output 	stream_address_17;
output 	stream_address_18;
output 	stream_address_19;
output 	stream_address_20;
output 	stream_address_21;
output 	stream_address_22;
output 	stream_address_23;
output 	stream_address_24;
output 	stream_address_25;
output 	stream_address_26;
output 	stream_address_27;
output 	stream_address_28;
output 	stream_address_29;
output 	stream_address_30;
output 	stream_address_31;
output 	user_reconfig_readdata_0;
input 	Equal3;
input 	basic_reconfig_readdata_0;
output 	user_reconfig_readdata_1;
input 	basic_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
input 	basic_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
input 	basic_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
input 	basic_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
output 	user_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
output 	user_reconfig_readdata_7;
input 	reconfig_mgmt_readdata_8;
input 	basic_reconfig_readdata_8;
output 	user_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
output 	user_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	user_reconfig_readdata_11;
output 	master_write;
input 	grant_7;
output 	mutex_req;
output 	mutex_grant;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
output 	stream_read;
output 	uif_busy;
input 	pll_mif_busy;
input 	ifsel_notdone_resync;
output 	uif_logical_ch_addr_0;
input 	comb;
output 	uif_logical_ch_addr_1;
output 	uif_logical_ch_addr_2;
output 	uif_logical_ch_addr_3;
input 	user_reconfig_readdata_101;
output 	uif_logical_ch_addr_4;
output 	uif_logical_ch_addr_5;
output 	uif_logical_ch_addr_6;
output 	uif_logical_ch_addr_7;
output 	uif_logical_ch_addr_8;
output 	uif_logical_ch_addr_9;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
output 	pll_go;
input 	uif_mode_0;
input 	Mux0;
input 	Mux3;
input 	WideOr0;
output 	pll_type;
output 	mif_rec_addr_7;
output 	mif_rec_addr_5;
output 	mif_rec_addr_6;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mif_waitrequest;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;
input 	reconfig_mif_readdata_15;
input 	reconfig_mif_readdata_14;
input 	reconfig_mif_readdata_13;
input 	reconfig_mif_readdata_12;
input 	reconfig_mif_readdata_11;
input 	reconfig_mif_readdata_1;
input 	reconfig_mif_readdata_0;
input 	reconfig_mif_readdata_4;
input 	reconfig_mif_readdata_3;
input 	reconfig_mif_readdata_2;
input 	reconfig_mif_readdata_7;
input 	reconfig_mif_readdata_5;
input 	reconfig_mif_readdata_6;
input 	reconfig_mif_readdata_8;
input 	reconfig_mif_readdata_9;
input 	reconfig_mif_readdata_10;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \inst_mif_ctrl|uif_rdata[5]~q ;
wire \inst_mif_ctrl|uif_rdata[6]~q ;
wire \inst_mif_ctrl|uif_rdata[7]~q ;
wire \inst_mif_ctrl|uif_rdata[8]~q ;
wire \inst_mif_ctrl|uif_rdata[9]~q ;
wire \inst_mif_ctrl|uif_rdata[10]~q ;
wire \inst_mif_ctrl|uif_rdata[11]~q ;
wire \inst_mif_ctrl|uif_rdata[12]~q ;
wire \inst_mif_ctrl|uif_rdata[13]~q ;
wire \inst_mif_ctrl|uif_rdata[14]~q ;
wire \inst_mif_ctrl|uif_rdata[15]~q ;
wire \inst_mif_ctrl|uif_rdata[16]~q ;
wire \inst_mif_ctrl|uif_rdata[17]~q ;
wire \inst_mif_ctrl|uif_rdata[18]~q ;
wire \inst_mif_ctrl|uif_rdata[19]~q ;
wire \inst_mif_ctrl|uif_rdata[20]~q ;
wire \inst_mif_ctrl|uif_rdata[21]~q ;
wire \inst_mif_ctrl|uif_rdata[22]~q ;
wire \inst_mif_ctrl|uif_rdata[23]~q ;
wire \inst_mif_ctrl|uif_rdata[24]~q ;
wire \inst_mif_ctrl|uif_rdata[25]~q ;
wire \inst_mif_ctrl|uif_rdata[26]~q ;
wire \inst_mif_ctrl|uif_rdata[27]~q ;
wire \inst_mif_ctrl|uif_rdata[28]~q ;
wire \inst_mif_ctrl|uif_rdata[29]~q ;
wire \inst_mif_ctrl|uif_rdata[30]~q ;
wire \inst_mif_ctrl|uif_rdata[31]~q ;
wire \inst_mif_ctrl|ctrl_addr[1]~q ;
wire \inst_mif_ctrl|ctrl_addr[2]~q ;
wire \inst_mif_ctrl|ctrl_addr[0]~q ;
wire \inst_mif_avmm|av_mif_addr[4]~q ;
wire \inst_mif_avmm|av_mif_addr[5]~q ;
wire \inst_mif_avmm|av_mif_addr[2]~q ;
wire \inst_mif_avmm|av_mif_addr[1]~q ;
wire \inst_mif_avmm|av_mif_addr[0]~q ;
wire \inst_mif_avmm|av_mif_addr[3]~q ;
wire \inst_mif_avmm|av_mif_addr[8]~q ;
wire \inst_mif_avmm|av_mif_addr[9]~q ;
wire \inst_mif_avmm|av_mif_addr[10]~q ;
wire \inst_mif_avmm|av_mif_addr[7]~q ;
wire \inst_mif_avmm|av_mif_addr[6]~q ;
wire \inst_mif_ctrl|ctrl_addr[4]~q ;
wire \inst_mif_ctrl|ctrl_addr[5]~q ;
wire \inst_mif_ctrl|ctrl_addr[6]~q ;
wire \inst_mif_ctrl|ctrl_addr[7]~q ;
wire \inst_mif_ctrl|ctrl_addr[8]~q ;
wire \inst_mif_ctrl|ctrl_addr[9]~q ;
wire \inst_mif_ctrl|ctrl_addr[10]~q ;
wire \inst_xreconf_uif|uif_writedata[0]~q ;
wire \inst_xreconf_uif|uif_mode[1]~q ;
wire \inst_xreconf_uif|uif_mode[0]~q ;
wire \inst_mif_ctrl|Equal5~0_combout ;
wire \inst_mif_ctrl|uif_rdata[0]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ;
wire \inst_xreconf_uif|uif_addr_offset[0]~q ;
wire \inst_xreconf_uif|uif_writedata[1]~q ;
wire \inst_mif_ctrl|uif_rdata[1]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ;
wire \inst_xreconf_uif|uif_addr_offset[1]~q ;
wire \inst_xreconf_uif|uif_writedata[2]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ;
wire \inst_xreconf_uif|uif_ctrl[0]~q ;
wire \inst_xreconf_uif|uif_addr_offset[2]~q ;
wire \inst_mif_ctrl|uif_rdata[2]~q ;
wire \inst_xreconf_uif|uif_writedata[3]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ;
wire \inst_xreconf_uif|uif_ctrl[1]~q ;
wire \inst_xreconf_uif|uif_addr_offset[3]~q ;
wire \inst_mif_ctrl|uif_rdata[3]~q ;
wire \inst_xreconf_uif|uif_writedata[4]~q ;
wire \inst_mif_ctrl|uif_rdata[4]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ;
wire \inst_xreconf_uif|uif_addr_offset[4]~q ;
wire \inst_xreconf_uif|uif_writedata[5]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ;
wire \inst_xreconf_uif|uif_addr_offset[5]~q ;
wire \inst_xreconf_uif|uif_writedata[6]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ;
wire \inst_xreconf_uif|uif_addr_offset[6]~q ;
wire \inst_xreconf_uif|uif_writedata[7]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ;
wire \inst_xreconf_uif|uif_addr_offset[7]~q ;
wire \inst_xreconf_uif|uif_writedata[8]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ;
wire \inst_xreconf_uif|uif_addr_offset[8]~q ;
wire \inst_xreconf_uif|uif_writedata[9]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ;
wire \inst_mif_ctrl|uif_addr_err~q ;
wire \inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ;
wire \inst_xreconf_uif|uif_addr_offset[9]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ;
wire \inst_xreconf_uif|uif_writedata[10]~q ;
wire \inst_xreconf_uif|uif_addr_offset[10]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ;
wire \inst_xreconf_uif|uif_writedata[11]~q ;
wire \inst_xreconf_uif|uif_addr_offset[11]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ;
wire \inst_xreconf_uif|uif_writedata[12]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ;
wire \inst_xreconf_uif|uif_writedata[13]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ;
wire \inst_xreconf_uif|uif_writedata[14]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ;
wire \inst_xreconf_uif|uif_writedata[15]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ;
wire \inst_xreconf_uif|uif_writedata[16]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ;
wire \inst_xreconf_uif|uif_writedata[17]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ;
wire \inst_xreconf_uif|uif_writedata[18]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ;
wire \inst_xreconf_uif|uif_writedata[19]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ;
wire \inst_xreconf_uif|uif_writedata[20]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ;
wire \inst_xreconf_uif|uif_writedata[21]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ;
wire \inst_xreconf_uif|uif_writedata[22]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ;
wire \inst_xreconf_uif|uif_writedata[23]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ;
wire \inst_xreconf_uif|uif_writedata[24]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ;
wire \inst_xreconf_uif|uif_writedata[25]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ;
wire \inst_xreconf_uif|uif_writedata[26]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ;
wire \inst_xreconf_uif|uif_writedata[27]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ;
wire \inst_xreconf_uif|uif_writedata[28]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ;
wire \inst_xreconf_uif|uif_writedata[29]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ;
wire \inst_xreconf_uif|uif_writedata[30]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ;
wire \inst_xreconf_uif|uif_writedata[31]~q ;
wire \inst_mif_ctrl|ctrl_opcode[1]~q ;
wire \inst_mif_ctrl|ctrl_opcode[2]~q ;
wire \inst_mif_ctrl|ctrl_opcode[0]~q ;
wire \inst_mif_ctrl|ctrl_go~q ;
wire \inst_mif_ctrl|ctrl_lock~q ;
wire \inst_mif_avmm|av_ctrl_req~q ;
wire \inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ;
wire \inst_mif_ctrl|ctrl_op_done~0_combout ;
wire \inst_mif_ctrl|mif_err_reg[4]~q ;
wire \inst_mif_ctrl|mif_err_reg[1]~q ;
wire \inst_mif_ctrl|mif_err_reg[0]~q ;
wire \inst_mif_ctrl|ctrl_av_go~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q ;
wire \inst_xreconf_uif|uif_go~q ;
wire \inst_mif_ctrl|mif_base_addr[0]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ;
wire \inst_mif_ctrl|mif_base_addr[1]~q ;
wire \inst_mif_ctrl|mif_base_addr[2]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ;
wire \inst_mif_ctrl|mif_base_addr[3]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ;
wire \inst_mif_ctrl|mif_base_addr[4]~q ;
wire \inst_mif_ctrl|mif_base_addr[5]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ;
wire \inst_mif_ctrl|mif_base_addr[6]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ;
wire \inst_mif_ctrl|mif_base_addr[7]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ;
wire \inst_mif_ctrl|mif_base_addr[8]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ;
wire \inst_mif_ctrl|mif_base_addr[9]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ;
wire \inst_mif_ctrl|mif_base_addr[10]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ;
wire \inst_mif_ctrl|mif_base_addr[11]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ;
wire \inst_mif_ctrl|mif_base_addr[12]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ;
wire \inst_mif_ctrl|mif_base_addr[13]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ;
wire \inst_mif_ctrl|mif_base_addr[14]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ;
wire \inst_mif_ctrl|mif_base_addr[15]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ;
wire \inst_mif_ctrl|mif_base_addr[16]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ;
wire \inst_mif_ctrl|mif_base_addr[17]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ;
wire \inst_mif_ctrl|mif_base_addr[18]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ;
wire \inst_mif_ctrl|mif_base_addr[19]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ;
wire \inst_mif_ctrl|mif_base_addr[20]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ;
wire \inst_mif_ctrl|mif_base_addr[21]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ;
wire \inst_mif_ctrl|mif_base_addr[22]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ;
wire \inst_mif_ctrl|mif_base_addr[23]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ;
wire \inst_mif_ctrl|mif_base_addr[24]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ;
wire \inst_mif_ctrl|mif_base_addr[25]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ;
wire \inst_mif_ctrl|mif_base_addr[26]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ;
wire \inst_mif_ctrl|mif_base_addr[27]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ;
wire \inst_mif_ctrl|mif_base_addr[28]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ;
wire \inst_mif_ctrl|mif_base_addr[29]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ;
wire \inst_mif_ctrl|mif_base_addr[30]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ;
wire \inst_mif_ctrl|mif_base_addr[31]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ;
wire \inst_mif_avmm|av_addr_burst~q ;
wire \inst_mif_ctrl|ctrl_wdata[1]~q ;
wire \inst_mif_ctrl|ctrl_wdata[2]~q ;
wire \inst_mif_ctrl|ctrl_wdata[0]~q ;
wire \inst_mif_ctrl|ctrl_wdata[3]~q ;
wire \inst_mif_ctrl|ctrl_addr[3]~q ;
wire \inst_mif_avmm|av_opcode_err~q ;
wire \inst_mif_ctrl|ctrl_wdata[4]~q ;
wire \inst_mif_ctrl|ctrl_wdata[5]~q ;
wire \inst_mif_ctrl|ctrl_wdata[6]~q ;
wire \inst_mif_ctrl|ctrl_wdata[7]~q ;
wire \inst_mif_ctrl|ctrl_wdata[8]~q ;
wire \inst_mif_ctrl|ctrl_wdata[9]~q ;
wire \inst_mif_ctrl|ctrl_wdata[10]~q ;
wire \inst_mif_ctrl|ctrl_wdata[11]~q ;
wire \inst_mif_ctrl|ctrl_addr[11]~q ;
wire \inst_mif_ctrl|ctrl_wdata[12]~q ;
wire \inst_mif_ctrl|ctrl_wdata[13]~q ;
wire \inst_mif_ctrl|ctrl_wdata[14]~q ;
wire \inst_mif_ctrl|ctrl_wdata[15]~q ;
wire \inst_mif_avmm|av_done~q ;
wire \inst_mif_avmm|mif_rec_data[1]~q ;
wire \inst_mif_avmm|mif_rec_data[2]~q ;
wire \inst_mif_avmm|mif_rec_data[0]~q ;
wire \inst_mif_avmm|mif_rec_data[3]~q ;
wire \inst_mif_avmm|av_mif_type_valid~q ;
wire \inst_mif_avmm|av_mif_type[1]~q ;
wire \inst_mif_avmm|av_mif_type[0]~q ;
wire \inst_mif_avmm|mif_rec_data[4]~q ;
wire \inst_mif_avmm|mif_rec_data[5]~q ;
wire \inst_mif_avmm|mif_rec_data[6]~q ;
wire \inst_mif_avmm|mif_rec_data[7]~q ;
wire \inst_mif_avmm|mif_rec_data[8]~q ;
wire \inst_mif_avmm|mif_rec_data[9]~q ;
wire \inst_mif_avmm|mif_rec_data[10]~q ;
wire \inst_mif_avmm|mif_rec_data[11]~q ;
wire \inst_mif_avmm|mif_rec_data[12]~q ;
wire \inst_mif_avmm|mif_rec_data[13]~q ;
wire \inst_mif_avmm|mif_rec_data[14]~q ;
wire \inst_mif_avmm|mif_rec_data[15]~q ;
wire \inst_mif_ctrl|mif_addr_mode~q ;


RECONFIGURE_IP_av_xcvr_reconfig_mif_ctrl inst_mif_ctrl(
	.uif_rdata_5(\inst_mif_ctrl|uif_rdata[5]~q ),
	.uif_rdata_6(\inst_mif_ctrl|uif_rdata[6]~q ),
	.uif_rdata_7(\inst_mif_ctrl|uif_rdata[7]~q ),
	.uif_rdata_8(\inst_mif_ctrl|uif_rdata[8]~q ),
	.uif_rdata_9(\inst_mif_ctrl|uif_rdata[9]~q ),
	.uif_rdata_10(\inst_mif_ctrl|uif_rdata[10]~q ),
	.uif_rdata_11(\inst_mif_ctrl|uif_rdata[11]~q ),
	.uif_rdata_12(\inst_mif_ctrl|uif_rdata[12]~q ),
	.uif_rdata_13(\inst_mif_ctrl|uif_rdata[13]~q ),
	.uif_rdata_14(\inst_mif_ctrl|uif_rdata[14]~q ),
	.uif_rdata_15(\inst_mif_ctrl|uif_rdata[15]~q ),
	.uif_rdata_16(\inst_mif_ctrl|uif_rdata[16]~q ),
	.uif_rdata_17(\inst_mif_ctrl|uif_rdata[17]~q ),
	.uif_rdata_18(\inst_mif_ctrl|uif_rdata[18]~q ),
	.uif_rdata_19(\inst_mif_ctrl|uif_rdata[19]~q ),
	.uif_rdata_20(\inst_mif_ctrl|uif_rdata[20]~q ),
	.uif_rdata_21(\inst_mif_ctrl|uif_rdata[21]~q ),
	.uif_rdata_22(\inst_mif_ctrl|uif_rdata[22]~q ),
	.uif_rdata_23(\inst_mif_ctrl|uif_rdata[23]~q ),
	.uif_rdata_24(\inst_mif_ctrl|uif_rdata[24]~q ),
	.uif_rdata_25(\inst_mif_ctrl|uif_rdata[25]~q ),
	.uif_rdata_26(\inst_mif_ctrl|uif_rdata[26]~q ),
	.uif_rdata_27(\inst_mif_ctrl|uif_rdata[27]~q ),
	.uif_rdata_28(\inst_mif_ctrl|uif_rdata[28]~q ),
	.uif_rdata_29(\inst_mif_ctrl|uif_rdata[29]~q ),
	.uif_rdata_30(\inst_mif_ctrl|uif_rdata[30]~q ),
	.uif_rdata_31(\inst_mif_ctrl|uif_rdata[31]~q ),
	.ctrl_addr_1(\inst_mif_ctrl|ctrl_addr[1]~q ),
	.ctrl_addr_2(\inst_mif_ctrl|ctrl_addr[2]~q ),
	.ctrl_addr_0(\inst_mif_ctrl|ctrl_addr[0]~q ),
	.av_mif_addr_4(\inst_mif_avmm|av_mif_addr[4]~q ),
	.av_mif_addr_5(\inst_mif_avmm|av_mif_addr[5]~q ),
	.av_mif_addr_2(\inst_mif_avmm|av_mif_addr[2]~q ),
	.av_mif_addr_1(\inst_mif_avmm|av_mif_addr[1]~q ),
	.av_mif_addr_0(\inst_mif_avmm|av_mif_addr[0]~q ),
	.av_mif_addr_3(\inst_mif_avmm|av_mif_addr[3]~q ),
	.av_mif_addr_8(\inst_mif_avmm|av_mif_addr[8]~q ),
	.av_mif_addr_9(\inst_mif_avmm|av_mif_addr[9]~q ),
	.av_mif_addr_10(\inst_mif_avmm|av_mif_addr[10]~q ),
	.av_mif_addr_7(\inst_mif_avmm|av_mif_addr[7]~q ),
	.av_mif_addr_6(\inst_mif_avmm|av_mif_addr[6]~q ),
	.ctrl_addr_4(\inst_mif_ctrl|ctrl_addr[4]~q ),
	.ctrl_addr_5(\inst_mif_ctrl|ctrl_addr[5]~q ),
	.ctrl_addr_6(\inst_mif_ctrl|ctrl_addr[6]~q ),
	.ctrl_addr_7(\inst_mif_ctrl|ctrl_addr[7]~q ),
	.ctrl_addr_8(\inst_mif_ctrl|ctrl_addr[8]~q ),
	.ctrl_addr_9(\inst_mif_ctrl|ctrl_addr[9]~q ),
	.ctrl_addr_10(\inst_mif_ctrl|ctrl_addr[10]~q ),
	.uif_busy1(uif_busy),
	.reset(ifsel_notdone_resync),
	.uif_writedata_0(\inst_xreconf_uif|uif_writedata[0]~q ),
	.uif_mode_1(\inst_xreconf_uif|uif_mode[1]~q ),
	.uif_mode_0(\inst_xreconf_uif|uif_mode[0]~q ),
	.Equal5(\inst_mif_ctrl|Equal5~0_combout ),
	.uif_rdata_0(\inst_mif_ctrl|uif_rdata[0]~q ),
	.uif_addr_offset_0(\inst_xreconf_uif|uif_addr_offset[0]~q ),
	.uif_writedata_1(\inst_xreconf_uif|uif_writedata[1]~q ),
	.uif_rdata_1(\inst_mif_ctrl|uif_rdata[1]~q ),
	.uif_addr_offset_1(\inst_xreconf_uif|uif_addr_offset[1]~q ),
	.uif_writedata_2(\inst_xreconf_uif|uif_writedata[2]~q ),
	.uif_ctrl_0(\inst_xreconf_uif|uif_ctrl[0]~q ),
	.uif_addr_offset_2(\inst_xreconf_uif|uif_addr_offset[2]~q ),
	.uif_rdata_2(\inst_mif_ctrl|uif_rdata[2]~q ),
	.uif_writedata_3(\inst_xreconf_uif|uif_writedata[3]~q ),
	.uif_ctrl_1(\inst_xreconf_uif|uif_ctrl[1]~q ),
	.uif_addr_offset_3(\inst_xreconf_uif|uif_addr_offset[3]~q ),
	.uif_rdata_3(\inst_mif_ctrl|uif_rdata[3]~q ),
	.uif_writedata_4(\inst_xreconf_uif|uif_writedata[4]~q ),
	.uif_rdata_4(\inst_mif_ctrl|uif_rdata[4]~q ),
	.uif_addr_offset_4(\inst_xreconf_uif|uif_addr_offset[4]~q ),
	.uif_writedata_5(\inst_xreconf_uif|uif_writedata[5]~q ),
	.uif_addr_offset_5(\inst_xreconf_uif|uif_addr_offset[5]~q ),
	.uif_writedata_6(\inst_xreconf_uif|uif_writedata[6]~q ),
	.uif_addr_offset_6(\inst_xreconf_uif|uif_addr_offset[6]~q ),
	.uif_writedata_7(\inst_xreconf_uif|uif_writedata[7]~q ),
	.uif_addr_offset_7(\inst_xreconf_uif|uif_addr_offset[7]~q ),
	.uif_writedata_8(\inst_xreconf_uif|uif_writedata[8]~q ),
	.uif_addr_offset_8(\inst_xreconf_uif|uif_addr_offset[8]~q ),
	.uif_writedata_9(\inst_xreconf_uif|uif_writedata[9]~q ),
	.uif_addr_err1(\inst_mif_ctrl|uif_addr_err~q ),
	.uif_addr_offset_9(\inst_xreconf_uif|uif_addr_offset[9]~q ),
	.uif_writedata_10(\inst_xreconf_uif|uif_writedata[10]~q ),
	.uif_addr_offset_10(\inst_xreconf_uif|uif_addr_offset[10]~q ),
	.uif_writedata_11(\inst_xreconf_uif|uif_writedata[11]~q ),
	.uif_addr_offset_11(\inst_xreconf_uif|uif_addr_offset[11]~q ),
	.uif_writedata_12(\inst_xreconf_uif|uif_writedata[12]~q ),
	.uif_writedata_13(\inst_xreconf_uif|uif_writedata[13]~q ),
	.uif_writedata_14(\inst_xreconf_uif|uif_writedata[14]~q ),
	.uif_writedata_15(\inst_xreconf_uif|uif_writedata[15]~q ),
	.uif_writedata_16(\inst_xreconf_uif|uif_writedata[16]~q ),
	.uif_writedata_17(\inst_xreconf_uif|uif_writedata[17]~q ),
	.uif_writedata_18(\inst_xreconf_uif|uif_writedata[18]~q ),
	.uif_writedata_19(\inst_xreconf_uif|uif_writedata[19]~q ),
	.uif_writedata_20(\inst_xreconf_uif|uif_writedata[20]~q ),
	.uif_writedata_21(\inst_xreconf_uif|uif_writedata[21]~q ),
	.uif_writedata_22(\inst_xreconf_uif|uif_writedata[22]~q ),
	.uif_writedata_23(\inst_xreconf_uif|uif_writedata[23]~q ),
	.uif_writedata_24(\inst_xreconf_uif|uif_writedata[24]~q ),
	.uif_writedata_25(\inst_xreconf_uif|uif_writedata[25]~q ),
	.uif_writedata_26(\inst_xreconf_uif|uif_writedata[26]~q ),
	.uif_writedata_27(\inst_xreconf_uif|uif_writedata[27]~q ),
	.uif_writedata_28(\inst_xreconf_uif|uif_writedata[28]~q ),
	.uif_writedata_29(\inst_xreconf_uif|uif_writedata[29]~q ),
	.uif_writedata_30(\inst_xreconf_uif|uif_writedata[30]~q ),
	.uif_writedata_31(\inst_xreconf_uif|uif_writedata[31]~q ),
	.ctrl_opcode_1(\inst_mif_ctrl|ctrl_opcode[1]~q ),
	.ctrl_opcode_2(\inst_mif_ctrl|ctrl_opcode[2]~q ),
	.ctrl_opcode_0(\inst_mif_ctrl|ctrl_opcode[0]~q ),
	.ctrl_go1(\inst_mif_ctrl|ctrl_go~q ),
	.ctrl_lock1(\inst_mif_ctrl|ctrl_lock~q ),
	.av_ctrl_req(\inst_mif_avmm|av_ctrl_req~q ),
	.waitrequest_to_ctrl(\inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ),
	.ctrl_op_done(\inst_mif_ctrl|ctrl_op_done~0_combout ),
	.mif_err_reg_4(\inst_mif_ctrl|mif_err_reg[4]~q ),
	.mif_err_reg_1(\inst_mif_ctrl|mif_err_reg[1]~q ),
	.mif_err_reg_0(\inst_mif_ctrl|mif_err_reg[0]~q ),
	.ctrl_av_go1(\inst_mif_ctrl|ctrl_av_go~q ),
	.ctrl_rdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q }),
	.uif_go(\inst_xreconf_uif|uif_go~q ),
	.mif_base_addr_0(\inst_mif_ctrl|mif_base_addr[0]~q ),
	.mif_base_addr_1(\inst_mif_ctrl|mif_base_addr[1]~q ),
	.mif_base_addr_2(\inst_mif_ctrl|mif_base_addr[2]~q ),
	.mif_base_addr_3(\inst_mif_ctrl|mif_base_addr[3]~q ),
	.mif_base_addr_4(\inst_mif_ctrl|mif_base_addr[4]~q ),
	.mif_base_addr_5(\inst_mif_ctrl|mif_base_addr[5]~q ),
	.mif_base_addr_6(\inst_mif_ctrl|mif_base_addr[6]~q ),
	.mif_base_addr_7(\inst_mif_ctrl|mif_base_addr[7]~q ),
	.mif_base_addr_8(\inst_mif_ctrl|mif_base_addr[8]~q ),
	.mif_base_addr_9(\inst_mif_ctrl|mif_base_addr[9]~q ),
	.mif_base_addr_10(\inst_mif_ctrl|mif_base_addr[10]~q ),
	.mif_base_addr_11(\inst_mif_ctrl|mif_base_addr[11]~q ),
	.mif_base_addr_12(\inst_mif_ctrl|mif_base_addr[12]~q ),
	.mif_base_addr_13(\inst_mif_ctrl|mif_base_addr[13]~q ),
	.mif_base_addr_14(\inst_mif_ctrl|mif_base_addr[14]~q ),
	.mif_base_addr_15(\inst_mif_ctrl|mif_base_addr[15]~q ),
	.mif_base_addr_16(\inst_mif_ctrl|mif_base_addr[16]~q ),
	.readdata_for_user_16(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.mif_base_addr_17(\inst_mif_ctrl|mif_base_addr[17]~q ),
	.readdata_for_user_17(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.mif_base_addr_18(\inst_mif_ctrl|mif_base_addr[18]~q ),
	.readdata_for_user_18(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.mif_base_addr_19(\inst_mif_ctrl|mif_base_addr[19]~q ),
	.readdata_for_user_19(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.mif_base_addr_20(\inst_mif_ctrl|mif_base_addr[20]~q ),
	.readdata_for_user_20(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.mif_base_addr_21(\inst_mif_ctrl|mif_base_addr[21]~q ),
	.readdata_for_user_21(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.mif_base_addr_22(\inst_mif_ctrl|mif_base_addr[22]~q ),
	.readdata_for_user_22(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.mif_base_addr_23(\inst_mif_ctrl|mif_base_addr[23]~q ),
	.readdata_for_user_23(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.mif_base_addr_24(\inst_mif_ctrl|mif_base_addr[24]~q ),
	.readdata_for_user_24(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.mif_base_addr_25(\inst_mif_ctrl|mif_base_addr[25]~q ),
	.readdata_for_user_25(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ),
	.mif_base_addr_26(\inst_mif_ctrl|mif_base_addr[26]~q ),
	.readdata_for_user_26(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ),
	.mif_base_addr_27(\inst_mif_ctrl|mif_base_addr[27]~q ),
	.readdata_for_user_27(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ),
	.mif_base_addr_28(\inst_mif_ctrl|mif_base_addr[28]~q ),
	.readdata_for_user_28(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ),
	.mif_base_addr_29(\inst_mif_ctrl|mif_base_addr[29]~q ),
	.readdata_for_user_29(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ),
	.mif_base_addr_30(\inst_mif_ctrl|mif_base_addr[30]~q ),
	.readdata_for_user_30(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ),
	.mif_base_addr_31(\inst_mif_ctrl|mif_base_addr[31]~q ),
	.readdata_for_user_31(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ),
	.av_addr_burst(\inst_mif_avmm|av_addr_burst~q ),
	.ctrl_wdata_1(\inst_mif_ctrl|ctrl_wdata[1]~q ),
	.ctrl_wdata_2(\inst_mif_ctrl|ctrl_wdata[2]~q ),
	.ctrl_wdata_0(\inst_mif_ctrl|ctrl_wdata[0]~q ),
	.ctrl_wdata_3(\inst_mif_ctrl|ctrl_wdata[3]~q ),
	.ctrl_addr_3(\inst_mif_ctrl|ctrl_addr[3]~q ),
	.av_opcode_err(\inst_mif_avmm|av_opcode_err~q ),
	.ctrl_wdata_4(\inst_mif_ctrl|ctrl_wdata[4]~q ),
	.ctrl_wdata_5(\inst_mif_ctrl|ctrl_wdata[5]~q ),
	.ctrl_wdata_6(\inst_mif_ctrl|ctrl_wdata[6]~q ),
	.ctrl_wdata_7(\inst_mif_ctrl|ctrl_wdata[7]~q ),
	.ctrl_wdata_8(\inst_mif_ctrl|ctrl_wdata[8]~q ),
	.ctrl_wdata_9(\inst_mif_ctrl|ctrl_wdata[9]~q ),
	.ctrl_wdata_10(\inst_mif_ctrl|ctrl_wdata[10]~q ),
	.ctrl_wdata_11(\inst_mif_ctrl|ctrl_wdata[11]~q ),
	.ctrl_addr_11(\inst_mif_ctrl|ctrl_addr[11]~q ),
	.ctrl_wdata_12(\inst_mif_ctrl|ctrl_wdata[12]~q ),
	.ctrl_wdata_13(\inst_mif_ctrl|ctrl_wdata[13]~q ),
	.ctrl_wdata_14(\inst_mif_ctrl|ctrl_wdata[14]~q ),
	.ctrl_wdata_15(\inst_mif_ctrl|ctrl_wdata[15]~q ),
	.av_done(\inst_mif_avmm|av_done~q ),
	.mif_rec_data_1(\inst_mif_avmm|mif_rec_data[1]~q ),
	.mif_rec_data_2(\inst_mif_avmm|mif_rec_data[2]~q ),
	.mif_rec_data_0(\inst_mif_avmm|mif_rec_data[0]~q ),
	.mif_rec_data_3(\inst_mif_avmm|mif_rec_data[3]~q ),
	.av_mif_type_valid(\inst_mif_avmm|av_mif_type_valid~q ),
	.av_mif_type_1(\inst_mif_avmm|av_mif_type[1]~q ),
	.av_mif_type_0(\inst_mif_avmm|av_mif_type[0]~q ),
	.mif_rec_data_4(\inst_mif_avmm|mif_rec_data[4]~q ),
	.mif_rec_data_5(\inst_mif_avmm|mif_rec_data[5]~q ),
	.mif_rec_data_6(\inst_mif_avmm|mif_rec_data[6]~q ),
	.mif_rec_data_7(\inst_mif_avmm|mif_rec_data[7]~q ),
	.mif_rec_data_8(\inst_mif_avmm|mif_rec_data[8]~q ),
	.mif_rec_data_9(\inst_mif_avmm|mif_rec_data[9]~q ),
	.mif_rec_data_10(\inst_mif_avmm|mif_rec_data[10]~q ),
	.mif_rec_data_11(\inst_mif_avmm|mif_rec_data[11]~q ),
	.mif_rec_data_12(\inst_mif_avmm|mif_rec_data[12]~q ),
	.mif_rec_data_13(\inst_mif_avmm|mif_rec_data[13]~q ),
	.mif_rec_data_14(\inst_mif_avmm|mif_rec_data[14]~q ),
	.mif_rec_data_15(\inst_mif_avmm|mif_rec_data[15]~q ),
	.mif_addr_mode1(\inst_mif_ctrl|mif_addr_mode~q ),
	.clk(mgmt_clk_clk));

RECONFIGURE_IP_alt_xreconf_uif_1 inst_xreconf_uif(
	.user_reconfig_readdata_12(user_reconfig_readdata_12),
	.user_reconfig_readdata_13(user_reconfig_readdata_13),
	.user_reconfig_readdata_14(user_reconfig_readdata_14),
	.user_reconfig_readdata_15(user_reconfig_readdata_15),
	.user_reconfig_readdata_16(user_reconfig_readdata_16),
	.user_reconfig_readdata_17(user_reconfig_readdata_17),
	.user_reconfig_readdata_18(user_reconfig_readdata_18),
	.user_reconfig_readdata_19(user_reconfig_readdata_19),
	.user_reconfig_readdata_20(user_reconfig_readdata_20),
	.user_reconfig_readdata_21(user_reconfig_readdata_21),
	.user_reconfig_readdata_22(user_reconfig_readdata_22),
	.user_reconfig_readdata_23(user_reconfig_readdata_23),
	.user_reconfig_readdata_24(user_reconfig_readdata_24),
	.user_reconfig_readdata_25(user_reconfig_readdata_25),
	.user_reconfig_readdata_26(user_reconfig_readdata_26),
	.user_reconfig_readdata_27(user_reconfig_readdata_27),
	.user_reconfig_readdata_28(user_reconfig_readdata_28),
	.user_reconfig_readdata_29(user_reconfig_readdata_29),
	.user_reconfig_readdata_30(user_reconfig_readdata_30),
	.user_reconfig_readdata_31(user_reconfig_readdata_31),
	.uif_rdata_5(\inst_mif_ctrl|uif_rdata[5]~q ),
	.uif_rdata_6(\inst_mif_ctrl|uif_rdata[6]~q ),
	.uif_rdata_7(\inst_mif_ctrl|uif_rdata[7]~q ),
	.uif_rdata_8(\inst_mif_ctrl|uif_rdata[8]~q ),
	.uif_rdata_9(\inst_mif_ctrl|uif_rdata[9]~q ),
	.uif_rdata_10(\inst_mif_ctrl|uif_rdata[10]~q ),
	.uif_rdata_11(\inst_mif_ctrl|uif_rdata[11]~q ),
	.uif_rdata_12(\inst_mif_ctrl|uif_rdata[12]~q ),
	.uif_rdata_13(\inst_mif_ctrl|uif_rdata[13]~q ),
	.uif_rdata_14(\inst_mif_ctrl|uif_rdata[14]~q ),
	.uif_rdata_15(\inst_mif_ctrl|uif_rdata[15]~q ),
	.uif_rdata_16(\inst_mif_ctrl|uif_rdata[16]~q ),
	.uif_rdata_17(\inst_mif_ctrl|uif_rdata[17]~q ),
	.uif_rdata_18(\inst_mif_ctrl|uif_rdata[18]~q ),
	.uif_rdata_19(\inst_mif_ctrl|uif_rdata[19]~q ),
	.uif_rdata_20(\inst_mif_ctrl|uif_rdata[20]~q ),
	.uif_rdata_21(\inst_mif_ctrl|uif_rdata[21]~q ),
	.uif_rdata_22(\inst_mif_ctrl|uif_rdata[22]~q ),
	.uif_rdata_23(\inst_mif_ctrl|uif_rdata[23]~q ),
	.uif_rdata_24(\inst_mif_ctrl|uif_rdata[24]~q ),
	.uif_rdata_25(\inst_mif_ctrl|uif_rdata[25]~q ),
	.uif_rdata_26(\inst_mif_ctrl|uif_rdata[26]~q ),
	.uif_rdata_27(\inst_mif_ctrl|uif_rdata[27]~q ),
	.uif_rdata_28(\inst_mif_ctrl|uif_rdata[28]~q ),
	.uif_rdata_29(\inst_mif_ctrl|uif_rdata[29]~q ),
	.uif_rdata_30(\inst_mif_ctrl|uif_rdata[30]~q ),
	.uif_rdata_31(\inst_mif_ctrl|uif_rdata[31]~q ),
	.user_reconfig_readdata_0(user_reconfig_readdata_0),
	.Equal3(Equal3),
	.user_reconfig_readdata_1(user_reconfig_readdata_1),
	.user_reconfig_readdata_2(user_reconfig_readdata_2),
	.user_reconfig_readdata_3(user_reconfig_readdata_3),
	.user_reconfig_readdata_4(user_reconfig_readdata_4),
	.user_reconfig_readdata_5(user_reconfig_readdata_5),
	.user_reconfig_readdata_6(user_reconfig_readdata_6),
	.user_reconfig_readdata_7(user_reconfig_readdata_7),
	.reconfig_mgmt_readdata_8(reconfig_mgmt_readdata_8),
	.user_reconfig_readdata_8(user_reconfig_readdata_8),
	.user_reconfig_readdata_9(user_reconfig_readdata_9),
	.user_reconfig_readdata_10(user_reconfig_readdata_10),
	.user_reconfig_readdata_11(user_reconfig_readdata_11),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg(launch_reg),
	.wait_reg(wait_reg),
	.uif_busy(uif_busy),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.uif_writedata_0(\inst_xreconf_uif|uif_writedata[0]~q ),
	.uif_mode_1(\inst_xreconf_uif|uif_mode[1]~q ),
	.uif_mode_0(\inst_xreconf_uif|uif_mode[0]~q ),
	.Equal5(\inst_mif_ctrl|Equal5~0_combout ),
	.uif_rdata_0(\inst_mif_ctrl|uif_rdata[0]~q ),
	.ph_readdata_0(\inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ),
	.uif_logical_ch_addr_0(uif_logical_ch_addr_0),
	.uif_addr_offset_0(\inst_xreconf_uif|uif_addr_offset[0]~q ),
	.comb(comb),
	.uif_writedata_1(\inst_xreconf_uif|uif_writedata[1]~q ),
	.uif_rdata_1(\inst_mif_ctrl|uif_rdata[1]~q ),
	.ph_readdata_1(\inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ),
	.uif_logical_ch_addr_1(uif_logical_ch_addr_1),
	.uif_addr_offset_1(\inst_xreconf_uif|uif_addr_offset[1]~q ),
	.uif_writedata_2(\inst_xreconf_uif|uif_writedata[2]~q ),
	.uif_logical_ch_addr_2(uif_logical_ch_addr_2),
	.ph_readdata_2(\inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ),
	.uif_ctrl_0(\inst_xreconf_uif|uif_ctrl[0]~q ),
	.uif_addr_offset_2(\inst_xreconf_uif|uif_addr_offset[2]~q ),
	.uif_rdata_2(\inst_mif_ctrl|uif_rdata[2]~q ),
	.uif_writedata_3(\inst_xreconf_uif|uif_writedata[3]~q ),
	.uif_logical_ch_addr_3(uif_logical_ch_addr_3),
	.ph_readdata_3(\inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ),
	.uif_ctrl_1(\inst_xreconf_uif|uif_ctrl[1]~q ),
	.uif_addr_offset_3(\inst_xreconf_uif|uif_addr_offset[3]~q ),
	.uif_rdata_3(\inst_mif_ctrl|uif_rdata[3]~q ),
	.user_reconfig_readdata_101(user_reconfig_readdata_101),
	.uif_writedata_4(\inst_xreconf_uif|uif_writedata[4]~q ),
	.uif_rdata_4(\inst_mif_ctrl|uif_rdata[4]~q ),
	.ph_readdata_4(\inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ),
	.uif_logical_ch_addr_4(uif_logical_ch_addr_4),
	.uif_addr_offset_4(\inst_xreconf_uif|uif_addr_offset[4]~q ),
	.uif_writedata_5(\inst_xreconf_uif|uif_writedata[5]~q ),
	.ph_readdata_5(\inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ),
	.uif_logical_ch_addr_5(uif_logical_ch_addr_5),
	.uif_addr_offset_5(\inst_xreconf_uif|uif_addr_offset[5]~q ),
	.uif_writedata_6(\inst_xreconf_uif|uif_writedata[6]~q ),
	.ph_readdata_6(\inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ),
	.uif_logical_ch_addr_6(uif_logical_ch_addr_6),
	.uif_addr_offset_6(\inst_xreconf_uif|uif_addr_offset[6]~q ),
	.uif_writedata_7(\inst_xreconf_uif|uif_writedata[7]~q ),
	.ph_readdata_7(\inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ),
	.uif_logical_ch_addr_7(uif_logical_ch_addr_7),
	.uif_addr_offset_7(\inst_xreconf_uif|uif_addr_offset[7]~q ),
	.uif_writedata_8(\inst_xreconf_uif|uif_writedata[8]~q ),
	.uif_logical_ch_addr_8(uif_logical_ch_addr_8),
	.ph_readdata_8(\inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ),
	.uif_addr_offset_8(\inst_xreconf_uif|uif_addr_offset[8]~q ),
	.uif_writedata_9(\inst_xreconf_uif|uif_writedata[9]~q ),
	.uif_logical_ch_addr_9(uif_logical_ch_addr_9),
	.ph_readdata_9(\inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ),
	.uif_addr_err(\inst_mif_ctrl|uif_addr_err~q ),
	.illegal_phy_ch(\inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ),
	.uif_addr_offset_9(\inst_xreconf_uif|uif_addr_offset[9]~q ),
	.ph_readdata_10(\inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ),
	.uif_writedata_10(\inst_xreconf_uif|uif_writedata[10]~q ),
	.uif_addr_offset_10(\inst_xreconf_uif|uif_addr_offset[10]~q ),
	.ph_readdata_11(\inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ),
	.uif_writedata_11(\inst_xreconf_uif|uif_writedata[11]~q ),
	.uif_addr_offset_11(\inst_xreconf_uif|uif_addr_offset[11]~q ),
	.ph_readdata_12(\inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ),
	.uif_writedata_12(\inst_xreconf_uif|uif_writedata[12]~q ),
	.ph_readdata_13(\inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ),
	.uif_writedata_13(\inst_xreconf_uif|uif_writedata[13]~q ),
	.ph_readdata_14(\inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ),
	.uif_writedata_14(\inst_xreconf_uif|uif_writedata[14]~q ),
	.ph_readdata_15(\inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ),
	.uif_writedata_15(\inst_xreconf_uif|uif_writedata[15]~q ),
	.ph_readdata_16(\inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ),
	.uif_writedata_16(\inst_xreconf_uif|uif_writedata[16]~q ),
	.ph_readdata_17(\inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ),
	.uif_writedata_17(\inst_xreconf_uif|uif_writedata[17]~q ),
	.ph_readdata_18(\inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ),
	.uif_writedata_18(\inst_xreconf_uif|uif_writedata[18]~q ),
	.ph_readdata_19(\inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ),
	.uif_writedata_19(\inst_xreconf_uif|uif_writedata[19]~q ),
	.ph_readdata_20(\inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ),
	.uif_writedata_20(\inst_xreconf_uif|uif_writedata[20]~q ),
	.ph_readdata_21(\inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ),
	.uif_writedata_21(\inst_xreconf_uif|uif_writedata[21]~q ),
	.ph_readdata_22(\inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ),
	.uif_writedata_22(\inst_xreconf_uif|uif_writedata[22]~q ),
	.ph_readdata_23(\inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ),
	.uif_writedata_23(\inst_xreconf_uif|uif_writedata[23]~q ),
	.ph_readdata_24(\inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ),
	.uif_writedata_24(\inst_xreconf_uif|uif_writedata[24]~q ),
	.ph_readdata_25(\inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ),
	.uif_writedata_25(\inst_xreconf_uif|uif_writedata[25]~q ),
	.ph_readdata_26(\inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ),
	.uif_writedata_26(\inst_xreconf_uif|uif_writedata[26]~q ),
	.ph_readdata_27(\inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ),
	.uif_writedata_27(\inst_xreconf_uif|uif_writedata[27]~q ),
	.ph_readdata_28(\inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ),
	.uif_writedata_28(\inst_xreconf_uif|uif_writedata[28]~q ),
	.ph_readdata_29(\inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ),
	.uif_writedata_29(\inst_xreconf_uif|uif_writedata[29]~q ),
	.ph_readdata_30(\inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ),
	.uif_writedata_30(\inst_xreconf_uif|uif_writedata[30]~q ),
	.ph_readdata_31(\inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ),
	.uif_writedata_31(\inst_xreconf_uif|uif_writedata[31]~q ),
	.uif_mode_01(uif_mode_0),
	.Mux0(Mux0),
	.Mux3(Mux3),
	.uif_go1(\inst_xreconf_uif|uif_go~q ),
	.WideOr0(WideOr0),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15));

RECONFIGURE_IP_alt_xreconf_cif_1 inst_xreconf_cif(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.ctrl_addr_1(\inst_mif_ctrl|ctrl_addr[1]~q ),
	.ctrl_addr_2(\inst_mif_ctrl|ctrl_addr[2]~q ),
	.ctrl_addr_0(\inst_mif_ctrl|ctrl_addr[0]~q ),
	.ctrl_addr_4(\inst_mif_ctrl|ctrl_addr[4]~q ),
	.ctrl_addr_5(\inst_mif_ctrl|ctrl_addr[5]~q ),
	.ctrl_addr_6(\inst_mif_ctrl|ctrl_addr[6]~q ),
	.ctrl_addr_7(\inst_mif_ctrl|ctrl_addr[7]~q ),
	.ctrl_addr_8(\inst_mif_ctrl|ctrl_addr[8]~q ),
	.ctrl_addr_9(\inst_mif_ctrl|ctrl_addr[9]~q ),
	.ctrl_addr_10(\inst_mif_ctrl|ctrl_addr[10]~q ),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.master_write(master_write),
	.grant_7(grant_7),
	.mutex_req(mutex_req),
	.mutex_grant(mutex_grant),
	.master_address_2(master_address_2),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.ph_readdata_0(\inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ),
	.uif_logical_ch_addr_0(uif_logical_ch_addr_0),
	.ph_readdata_1(\inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ),
	.uif_logical_ch_addr_1(uif_logical_ch_addr_1),
	.uif_logical_ch_addr_2(uif_logical_ch_addr_2),
	.ph_readdata_2(\inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ),
	.uif_logical_ch_addr_3(uif_logical_ch_addr_3),
	.ph_readdata_3(\inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ),
	.ph_readdata_4(\inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ),
	.uif_logical_ch_addr_4(uif_logical_ch_addr_4),
	.ph_readdata_5(\inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ),
	.uif_logical_ch_addr_5(uif_logical_ch_addr_5),
	.ph_readdata_6(\inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ),
	.uif_logical_ch_addr_6(uif_logical_ch_addr_6),
	.ph_readdata_7(\inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ),
	.uif_logical_ch_addr_7(uif_logical_ch_addr_7),
	.uif_logical_ch_addr_8(uif_logical_ch_addr_8),
	.ph_readdata_8(\inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ),
	.uif_logical_ch_addr_9(uif_logical_ch_addr_9),
	.ph_readdata_9(\inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ),
	.illegal_phy_ch(\inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ),
	.ph_readdata_10(\inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ),
	.ph_readdata_11(\inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ),
	.ph_readdata_12(\inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ),
	.ph_readdata_13(\inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ),
	.ph_readdata_14(\inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ),
	.ph_readdata_15(\inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ),
	.ph_readdata_16(\inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ),
	.ph_readdata_17(\inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ),
	.ph_readdata_18(\inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ),
	.ph_readdata_19(\inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ),
	.ph_readdata_20(\inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ),
	.ph_readdata_21(\inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ),
	.ph_readdata_22(\inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ),
	.ph_readdata_23(\inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ),
	.ph_readdata_24(\inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ),
	.ph_readdata_25(\inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ),
	.ph_readdata_26(\inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ),
	.ph_readdata_27(\inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ),
	.ph_readdata_28(\inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ),
	.ph_readdata_29(\inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ),
	.ph_readdata_30(\inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ),
	.ph_readdata_31(\inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.ctrl_opcode_1(\inst_mif_ctrl|ctrl_opcode[1]~q ),
	.ctrl_opcode_2(\inst_mif_ctrl|ctrl_opcode[2]~q ),
	.ctrl_opcode_0(\inst_mif_ctrl|ctrl_opcode[0]~q ),
	.ctrl_go(\inst_mif_ctrl|ctrl_go~q ),
	.ctrl_lock(\inst_mif_ctrl|ctrl_lock~q ),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.waitrequest_to_ctrl(\inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.master_writedata_11(master_writedata_11),
	.master_writedata_12(master_writedata_12),
	.master_writedata_13(master_writedata_13),
	.master_writedata_14(master_writedata_14),
	.master_writedata_15(master_writedata_15),
	.readdata_for_user_0(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q ),
	.readdata_for_user_1(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ),
	.readdata_for_user_2(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ),
	.readdata_for_user_3(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ),
	.readdata_for_user_4(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ),
	.readdata_for_user_5(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ),
	.readdata_for_user_6(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ),
	.readdata_for_user_7(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ),
	.readdata_for_user_8(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ),
	.readdata_for_user_9(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ),
	.readdata_for_user_10(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ),
	.readdata_for_user_11(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ),
	.readdata_for_user_12(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ),
	.readdata_for_user_13(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ),
	.readdata_for_user_14(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ),
	.readdata_for_user_15(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ),
	.readdata_for_user_16(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.readdata_for_user_17(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.readdata_for_user_18(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.readdata_for_user_19(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.readdata_for_user_20(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.readdata_for_user_21(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.readdata_for_user_22(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.readdata_for_user_23(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.readdata_for_user_24(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.readdata_for_user_25(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[25]~q ),
	.readdata_for_user_26(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[26]~q ),
	.readdata_for_user_27(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[27]~q ),
	.readdata_for_user_28(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[28]~q ),
	.readdata_for_user_29(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[29]~q ),
	.readdata_for_user_30(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[30]~q ),
	.readdata_for_user_31(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[31]~q ),
	.ctrl_wdata_1(\inst_mif_ctrl|ctrl_wdata[1]~q ),
	.ctrl_wdata_2(\inst_mif_ctrl|ctrl_wdata[2]~q ),
	.ctrl_wdata_0(\inst_mif_ctrl|ctrl_wdata[0]~q ),
	.ctrl_wdata_3(\inst_mif_ctrl|ctrl_wdata[3]~q ),
	.ctrl_addr_3(\inst_mif_ctrl|ctrl_addr[3]~q ),
	.ctrl_wdata_4(\inst_mif_ctrl|ctrl_wdata[4]~q ),
	.ctrl_wdata_5(\inst_mif_ctrl|ctrl_wdata[5]~q ),
	.ctrl_wdata_6(\inst_mif_ctrl|ctrl_wdata[6]~q ),
	.ctrl_wdata_7(\inst_mif_ctrl|ctrl_wdata[7]~q ),
	.ctrl_wdata_8(\inst_mif_ctrl|ctrl_wdata[8]~q ),
	.ctrl_wdata_9(\inst_mif_ctrl|ctrl_wdata[9]~q ),
	.ctrl_wdata_10(\inst_mif_ctrl|ctrl_wdata[10]~q ),
	.ctrl_wdata_11(\inst_mif_ctrl|ctrl_wdata[11]~q ),
	.ctrl_addr_11(\inst_mif_ctrl|ctrl_addr[11]~q ),
	.ctrl_wdata_12(\inst_mif_ctrl|ctrl_wdata[12]~q ),
	.ctrl_wdata_13(\inst_mif_ctrl|ctrl_wdata[13]~q ),
	.ctrl_wdata_14(\inst_mif_ctrl|ctrl_wdata[14]~q ),
	.ctrl_wdata_15(\inst_mif_ctrl|ctrl_wdata[15]~q ),
	.mgmt_clk_clk(mgmt_clk_clk));

RECONFIGURE_IP_av_xcvr_reconfig_mif_avmm inst_mif_avmm(
	.stream_address_0(stream_address_0),
	.stream_address_1(stream_address_1),
	.stream_address_2(stream_address_2),
	.stream_address_3(stream_address_3),
	.stream_address_4(stream_address_4),
	.stream_address_5(stream_address_5),
	.stream_address_6(stream_address_6),
	.stream_address_7(stream_address_7),
	.stream_address_8(stream_address_8),
	.stream_address_9(stream_address_9),
	.stream_address_10(stream_address_10),
	.stream_address_11(stream_address_11),
	.stream_address_12(stream_address_12),
	.stream_address_13(stream_address_13),
	.stream_address_14(stream_address_14),
	.stream_address_15(stream_address_15),
	.stream_address_16(stream_address_16),
	.stream_address_17(stream_address_17),
	.stream_address_18(stream_address_18),
	.stream_address_19(stream_address_19),
	.stream_address_20(stream_address_20),
	.stream_address_21(stream_address_21),
	.stream_address_22(stream_address_22),
	.stream_address_23(stream_address_23),
	.stream_address_24(stream_address_24),
	.stream_address_25(stream_address_25),
	.stream_address_26(stream_address_26),
	.stream_address_27(stream_address_27),
	.stream_address_28(stream_address_28),
	.stream_address_29(stream_address_29),
	.stream_address_30(stream_address_30),
	.stream_address_31(stream_address_31),
	.av_mif_addr_4(\inst_mif_avmm|av_mif_addr[4]~q ),
	.av_mif_addr_5(\inst_mif_avmm|av_mif_addr[5]~q ),
	.av_mif_addr_2(\inst_mif_avmm|av_mif_addr[2]~q ),
	.av_mif_addr_1(\inst_mif_avmm|av_mif_addr[1]~q ),
	.av_mif_addr_0(\inst_mif_avmm|av_mif_addr[0]~q ),
	.av_mif_addr_3(\inst_mif_avmm|av_mif_addr[3]~q ),
	.av_mif_addr_8(\inst_mif_avmm|av_mif_addr[8]~q ),
	.av_mif_addr_9(\inst_mif_avmm|av_mif_addr[9]~q ),
	.av_mif_addr_10(\inst_mif_avmm|av_mif_addr[10]~q ),
	.av_mif_addr_7(\inst_mif_avmm|av_mif_addr[7]~q ),
	.av_mif_addr_6(\inst_mif_avmm|av_mif_addr[6]~q ),
	.stream_read1(stream_read),
	.pll_mif_busy(pll_mif_busy),
	.reset(ifsel_notdone_resync),
	.av_ctrl_req1(\inst_mif_avmm|av_ctrl_req~q ),
	.ctrl_op_done(\inst_mif_ctrl|ctrl_op_done~0_combout ),
	.mif_err_reg_4(\inst_mif_ctrl|mif_err_reg[4]~q ),
	.mif_err_reg_1(\inst_mif_ctrl|mif_err_reg[1]~q ),
	.mif_err_reg_0(\inst_mif_ctrl|mif_err_reg[0]~q ),
	.ctrl_av_go(\inst_mif_ctrl|ctrl_av_go~q ),
	.pll_go1(pll_go),
	.mif_base_addr_0(\inst_mif_ctrl|mif_base_addr[0]~q ),
	.mif_base_addr_1(\inst_mif_ctrl|mif_base_addr[1]~q ),
	.mif_base_addr_2(\inst_mif_ctrl|mif_base_addr[2]~q ),
	.mif_base_addr_3(\inst_mif_ctrl|mif_base_addr[3]~q ),
	.mif_base_addr_4(\inst_mif_ctrl|mif_base_addr[4]~q ),
	.mif_base_addr_5(\inst_mif_ctrl|mif_base_addr[5]~q ),
	.mif_base_addr_6(\inst_mif_ctrl|mif_base_addr[6]~q ),
	.mif_base_addr_7(\inst_mif_ctrl|mif_base_addr[7]~q ),
	.mif_base_addr_8(\inst_mif_ctrl|mif_base_addr[8]~q ),
	.mif_base_addr_9(\inst_mif_ctrl|mif_base_addr[9]~q ),
	.mif_base_addr_10(\inst_mif_ctrl|mif_base_addr[10]~q ),
	.mif_base_addr_11(\inst_mif_ctrl|mif_base_addr[11]~q ),
	.mif_base_addr_12(\inst_mif_ctrl|mif_base_addr[12]~q ),
	.mif_base_addr_13(\inst_mif_ctrl|mif_base_addr[13]~q ),
	.mif_base_addr_14(\inst_mif_ctrl|mif_base_addr[14]~q ),
	.mif_base_addr_15(\inst_mif_ctrl|mif_base_addr[15]~q ),
	.mif_base_addr_16(\inst_mif_ctrl|mif_base_addr[16]~q ),
	.mif_base_addr_17(\inst_mif_ctrl|mif_base_addr[17]~q ),
	.mif_base_addr_18(\inst_mif_ctrl|mif_base_addr[18]~q ),
	.mif_base_addr_19(\inst_mif_ctrl|mif_base_addr[19]~q ),
	.mif_base_addr_20(\inst_mif_ctrl|mif_base_addr[20]~q ),
	.mif_base_addr_21(\inst_mif_ctrl|mif_base_addr[21]~q ),
	.mif_base_addr_22(\inst_mif_ctrl|mif_base_addr[22]~q ),
	.mif_base_addr_23(\inst_mif_ctrl|mif_base_addr[23]~q ),
	.mif_base_addr_24(\inst_mif_ctrl|mif_base_addr[24]~q ),
	.mif_base_addr_25(\inst_mif_ctrl|mif_base_addr[25]~q ),
	.mif_base_addr_26(\inst_mif_ctrl|mif_base_addr[26]~q ),
	.mif_base_addr_27(\inst_mif_ctrl|mif_base_addr[27]~q ),
	.mif_base_addr_28(\inst_mif_ctrl|mif_base_addr[28]~q ),
	.mif_base_addr_29(\inst_mif_ctrl|mif_base_addr[29]~q ),
	.mif_base_addr_30(\inst_mif_ctrl|mif_base_addr[30]~q ),
	.mif_base_addr_31(\inst_mif_ctrl|mif_base_addr[31]~q ),
	.av_addr_burst1(\inst_mif_avmm|av_addr_burst~q ),
	.av_opcode_err1(\inst_mif_avmm|av_opcode_err~q ),
	.av_done1(\inst_mif_avmm|av_done~q ),
	.pll_type1(pll_type),
	.mif_rec_data_1(\inst_mif_avmm|mif_rec_data[1]~q ),
	.mif_rec_addr_7(mif_rec_addr_7),
	.mif_rec_addr_5(mif_rec_addr_5),
	.mif_rec_addr_6(mif_rec_addr_6),
	.mif_rec_data_2(\inst_mif_avmm|mif_rec_data[2]~q ),
	.mif_rec_data_0(\inst_mif_avmm|mif_rec_data[0]~q ),
	.mif_rec_data_3(\inst_mif_avmm|mif_rec_data[3]~q ),
	.av_mif_type_valid1(\inst_mif_avmm|av_mif_type_valid~q ),
	.av_mif_type_1(\inst_mif_avmm|av_mif_type[1]~q ),
	.av_mif_type_0(\inst_mif_avmm|av_mif_type[0]~q ),
	.mif_rec_data_4(\inst_mif_avmm|mif_rec_data[4]~q ),
	.mif_rec_data_5(\inst_mif_avmm|mif_rec_data[5]~q ),
	.mif_rec_data_6(\inst_mif_avmm|mif_rec_data[6]~q ),
	.mif_rec_data_7(\inst_mif_avmm|mif_rec_data[7]~q ),
	.mif_rec_data_8(\inst_mif_avmm|mif_rec_data[8]~q ),
	.mif_rec_data_9(\inst_mif_avmm|mif_rec_data[9]~q ),
	.mif_rec_data_10(\inst_mif_avmm|mif_rec_data[10]~q ),
	.mif_rec_data_11(\inst_mif_avmm|mif_rec_data[11]~q ),
	.mif_rec_data_12(\inst_mif_avmm|mif_rec_data[12]~q ),
	.mif_rec_data_13(\inst_mif_avmm|mif_rec_data[13]~q ),
	.mif_rec_data_14(\inst_mif_avmm|mif_rec_data[14]~q ),
	.mif_rec_data_15(\inst_mif_avmm|mif_rec_data[15]~q ),
	.mif_addr_mode(\inst_mif_ctrl|mif_addr_mode~q ),
	.clk(mgmt_clk_clk),
	.reconfig_mif_waitrequest(reconfig_mif_waitrequest),
	.stream_readdata({reconfig_mif_readdata_15,reconfig_mif_readdata_14,reconfig_mif_readdata_13,reconfig_mif_readdata_12,reconfig_mif_readdata_11,reconfig_mif_readdata_10,reconfig_mif_readdata_9,reconfig_mif_readdata_8,reconfig_mif_readdata_7,reconfig_mif_readdata_6,
reconfig_mif_readdata_5,reconfig_mif_readdata_4,reconfig_mif_readdata_3,reconfig_mif_readdata_2,reconfig_mif_readdata_1,reconfig_mif_readdata_0}));

endmodule

module RECONFIGURE_IP_alt_xreconf_cif_1 (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	ctrl_addr_1,
	ctrl_addr_2,
	ctrl_addr_0,
	ctrl_addr_4,
	ctrl_addr_5,
	ctrl_addr_6,
	ctrl_addr_7,
	ctrl_addr_8,
	ctrl_addr_9,
	ctrl_addr_10,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write,
	grant_7,
	mutex_req,
	mutex_grant,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	ifsel_notdone_resync,
	ph_readdata_0,
	uif_logical_ch_addr_0,
	ph_readdata_1,
	uif_logical_ch_addr_1,
	uif_logical_ch_addr_2,
	ph_readdata_2,
	uif_logical_ch_addr_3,
	ph_readdata_3,
	ph_readdata_4,
	uif_logical_ch_addr_4,
	ph_readdata_5,
	uif_logical_ch_addr_5,
	ph_readdata_6,
	uif_logical_ch_addr_6,
	ph_readdata_7,
	uif_logical_ch_addr_7,
	uif_logical_ch_addr_8,
	ph_readdata_8,
	uif_logical_ch_addr_9,
	ph_readdata_9,
	illegal_phy_ch,
	ph_readdata_10,
	ph_readdata_11,
	ph_readdata_12,
	ph_readdata_13,
	ph_readdata_14,
	ph_readdata_15,
	ph_readdata_16,
	ph_readdata_17,
	ph_readdata_18,
	ph_readdata_19,
	ph_readdata_20,
	ph_readdata_21,
	ph_readdata_22,
	ph_readdata_23,
	ph_readdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	ctrl_opcode_1,
	ctrl_opcode_2,
	ctrl_opcode_0,
	ctrl_go,
	ctrl_lock,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	waitrequest_to_ctrl,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	readdata_for_user_0,
	readdata_for_user_1,
	readdata_for_user_2,
	readdata_for_user_3,
	readdata_for_user_4,
	readdata_for_user_5,
	readdata_for_user_6,
	readdata_for_user_7,
	readdata_for_user_8,
	readdata_for_user_9,
	readdata_for_user_10,
	readdata_for_user_11,
	readdata_for_user_12,
	readdata_for_user_13,
	readdata_for_user_14,
	readdata_for_user_15,
	readdata_for_user_16,
	readdata_for_user_17,
	readdata_for_user_18,
	readdata_for_user_19,
	readdata_for_user_20,
	readdata_for_user_21,
	readdata_for_user_22,
	readdata_for_user_23,
	readdata_for_user_24,
	readdata_for_user_25,
	readdata_for_user_26,
	readdata_for_user_27,
	readdata_for_user_28,
	readdata_for_user_29,
	readdata_for_user_30,
	readdata_for_user_31,
	ctrl_wdata_1,
	ctrl_wdata_2,
	ctrl_wdata_0,
	ctrl_wdata_3,
	ctrl_addr_3,
	ctrl_wdata_4,
	ctrl_wdata_5,
	ctrl_wdata_6,
	ctrl_wdata_7,
	ctrl_wdata_8,
	ctrl_wdata_9,
	ctrl_wdata_10,
	ctrl_wdata_11,
	ctrl_addr_11,
	ctrl_wdata_12,
	ctrl_wdata_13,
	ctrl_wdata_14,
	ctrl_wdata_15,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_16;
input 	basic_reconfig_readdata_17;
input 	basic_reconfig_readdata_18;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
input 	ctrl_addr_1;
input 	ctrl_addr_2;
input 	ctrl_addr_0;
input 	ctrl_addr_4;
input 	ctrl_addr_5;
input 	ctrl_addr_6;
input 	ctrl_addr_7;
input 	ctrl_addr_8;
input 	ctrl_addr_9;
input 	ctrl_addr_10;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write;
input 	grant_7;
output 	mutex_req;
output 	mutex_grant;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	ifsel_notdone_resync;
output 	ph_readdata_0;
input 	uif_logical_ch_addr_0;
output 	ph_readdata_1;
input 	uif_logical_ch_addr_1;
input 	uif_logical_ch_addr_2;
output 	ph_readdata_2;
input 	uif_logical_ch_addr_3;
output 	ph_readdata_3;
output 	ph_readdata_4;
input 	uif_logical_ch_addr_4;
output 	ph_readdata_5;
input 	uif_logical_ch_addr_5;
output 	ph_readdata_6;
input 	uif_logical_ch_addr_6;
output 	ph_readdata_7;
input 	uif_logical_ch_addr_7;
input 	uif_logical_ch_addr_8;
output 	ph_readdata_8;
input 	uif_logical_ch_addr_9;
output 	ph_readdata_9;
output 	illegal_phy_ch;
output 	ph_readdata_10;
output 	ph_readdata_11;
output 	ph_readdata_12;
output 	ph_readdata_13;
output 	ph_readdata_14;
output 	ph_readdata_15;
output 	ph_readdata_16;
output 	ph_readdata_17;
output 	ph_readdata_18;
output 	ph_readdata_19;
output 	ph_readdata_20;
output 	ph_readdata_21;
output 	ph_readdata_22;
output 	ph_readdata_23;
output 	ph_readdata_24;
output 	ph_readdata_25;
output 	ph_readdata_26;
output 	ph_readdata_27;
output 	ph_readdata_28;
output 	ph_readdata_29;
output 	ph_readdata_30;
output 	ph_readdata_31;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
input 	ctrl_opcode_1;
input 	ctrl_opcode_2;
input 	ctrl_opcode_0;
input 	ctrl_go;
input 	ctrl_lock;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	waitrequest_to_ctrl;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
output 	readdata_for_user_0;
output 	readdata_for_user_1;
output 	readdata_for_user_2;
output 	readdata_for_user_3;
output 	readdata_for_user_4;
output 	readdata_for_user_5;
output 	readdata_for_user_6;
output 	readdata_for_user_7;
output 	readdata_for_user_8;
output 	readdata_for_user_9;
output 	readdata_for_user_10;
output 	readdata_for_user_11;
output 	readdata_for_user_12;
output 	readdata_for_user_13;
output 	readdata_for_user_14;
output 	readdata_for_user_15;
output 	readdata_for_user_16;
output 	readdata_for_user_17;
output 	readdata_for_user_18;
output 	readdata_for_user_19;
output 	readdata_for_user_20;
output 	readdata_for_user_21;
output 	readdata_for_user_22;
output 	readdata_for_user_23;
output 	readdata_for_user_24;
output 	readdata_for_user_25;
output 	readdata_for_user_26;
output 	readdata_for_user_27;
output 	readdata_for_user_28;
output 	readdata_for_user_29;
output 	readdata_for_user_30;
output 	readdata_for_user_31;
input 	ctrl_wdata_1;
input 	ctrl_wdata_2;
input 	ctrl_wdata_0;
input 	ctrl_wdata_3;
input 	ctrl_addr_3;
input 	ctrl_wdata_4;
input 	ctrl_wdata_5;
input 	ctrl_wdata_6;
input 	ctrl_wdata_7;
input 	ctrl_wdata_8;
input 	ctrl_wdata_9;
input 	ctrl_wdata_10;
input 	ctrl_wdata_11;
input 	ctrl_addr_11;
input 	ctrl_wdata_12;
input 	ctrl_wdata_13;
input 	ctrl_wdata_14;
input 	ctrl_wdata_15;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



RECONFIGURE_IP_alt_arbiter_acq_2 mutex_inst(
	.grant_7(grant_7),
	.mutex_req(mutex_req),
	.mutex_grant1(mutex_grant));

RECONFIGURE_IP_alt_xreconf_basic_acq_1 inst_basic_acq(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.ctrl_addr_1(ctrl_addr_1),
	.ctrl_addr_2(ctrl_addr_2),
	.ctrl_addr_0(ctrl_addr_0),
	.ctrl_addr_4(ctrl_addr_4),
	.ctrl_addr_5(ctrl_addr_5),
	.ctrl_addr_6(ctrl_addr_6),
	.ctrl_addr_7(ctrl_addr_7),
	.ctrl_addr_8(ctrl_addr_8),
	.ctrl_addr_9(ctrl_addr_9),
	.ctrl_addr_10(ctrl_addr_10),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.master_write1(master_write),
	.mutex_req1(mutex_req),
	.mutex_grant(mutex_grant),
	.master_address_2(master_address_2),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read1(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.reset(ifsel_notdone_resync),
	.ph_readdata_0(ph_readdata_0),
	.logical_ch_addr({uif_logical_ch_addr_9,uif_logical_ch_addr_8,uif_logical_ch_addr_7,uif_logical_ch_addr_6,uif_logical_ch_addr_5,uif_logical_ch_addr_4,uif_logical_ch_addr_3,uif_logical_ch_addr_2,uif_logical_ch_addr_1,uif_logical_ch_addr_0}),
	.ph_readdata_1(ph_readdata_1),
	.ph_readdata_2(ph_readdata_2),
	.ph_readdata_3(ph_readdata_3),
	.ph_readdata_4(ph_readdata_4),
	.ph_readdata_5(ph_readdata_5),
	.ph_readdata_6(ph_readdata_6),
	.ph_readdata_7(ph_readdata_7),
	.ph_readdata_8(ph_readdata_8),
	.ph_readdata_9(ph_readdata_9),
	.illegal_phy_ch1(illegal_phy_ch),
	.ph_readdata_10(ph_readdata_10),
	.ph_readdata_11(ph_readdata_11),
	.ph_readdata_12(ph_readdata_12),
	.ph_readdata_13(ph_readdata_13),
	.ph_readdata_14(ph_readdata_14),
	.ph_readdata_15(ph_readdata_15),
	.ph_readdata_16(ph_readdata_16),
	.ph_readdata_17(ph_readdata_17),
	.ph_readdata_18(ph_readdata_18),
	.ph_readdata_19(ph_readdata_19),
	.ph_readdata_20(ph_readdata_20),
	.ph_readdata_21(ph_readdata_21),
	.ph_readdata_22(ph_readdata_22),
	.ph_readdata_23(ph_readdata_23),
	.ph_readdata_24(ph_readdata_24),
	.ph_readdata_25(ph_readdata_25),
	.ph_readdata_26(ph_readdata_26),
	.ph_readdata_27(ph_readdata_27),
	.ph_readdata_28(ph_readdata_28),
	.ph_readdata_29(ph_readdata_29),
	.ph_readdata_30(ph_readdata_30),
	.ph_readdata_31(ph_readdata_31),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.ctrl_opcode_1(ctrl_opcode_1),
	.ctrl_opcode_2(ctrl_opcode_2),
	.ctrl_opcode_0(ctrl_opcode_0),
	.ctrl_go(ctrl_go),
	.ctrl_lock(ctrl_lock),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.waitrequest_to_ctrl1(waitrequest_to_ctrl),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.master_writedata_11(master_writedata_11),
	.master_writedata_12(master_writedata_12),
	.master_writedata_13(master_writedata_13),
	.master_writedata_14(master_writedata_14),
	.master_writedata_15(master_writedata_15),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_1(readdata_for_user_1),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_9(readdata_for_user_9),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_13(readdata_for_user_13),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_16(readdata_for_user_16),
	.readdata_for_user_17(readdata_for_user_17),
	.readdata_for_user_18(readdata_for_user_18),
	.readdata_for_user_19(readdata_for_user_19),
	.readdata_for_user_20(readdata_for_user_20),
	.readdata_for_user_21(readdata_for_user_21),
	.readdata_for_user_22(readdata_for_user_22),
	.readdata_for_user_23(readdata_for_user_23),
	.readdata_for_user_24(readdata_for_user_24),
	.readdata_for_user_25(readdata_for_user_25),
	.readdata_for_user_26(readdata_for_user_26),
	.readdata_for_user_27(readdata_for_user_27),
	.readdata_for_user_28(readdata_for_user_28),
	.readdata_for_user_29(readdata_for_user_29),
	.readdata_for_user_30(readdata_for_user_30),
	.readdata_for_user_31(readdata_for_user_31),
	.ctrl_wdata_1(ctrl_wdata_1),
	.ctrl_wdata_2(ctrl_wdata_2),
	.ctrl_wdata_0(ctrl_wdata_0),
	.ctrl_wdata_3(ctrl_wdata_3),
	.ctrl_addr_3(ctrl_addr_3),
	.ctrl_wdata_4(ctrl_wdata_4),
	.ctrl_wdata_5(ctrl_wdata_5),
	.ctrl_wdata_6(ctrl_wdata_6),
	.ctrl_wdata_7(ctrl_wdata_7),
	.ctrl_wdata_8(ctrl_wdata_8),
	.ctrl_wdata_9(ctrl_wdata_9),
	.ctrl_wdata_10(ctrl_wdata_10),
	.ctrl_wdata_11(ctrl_wdata_11),
	.ctrl_addr_11(ctrl_addr_11),
	.ctrl_wdata_12(ctrl_wdata_12),
	.ctrl_wdata_13(ctrl_wdata_13),
	.ctrl_wdata_14(ctrl_wdata_14),
	.ctrl_wdata_15(ctrl_wdata_15),
	.clk(mgmt_clk_clk));

endmodule

module RECONFIGURE_IP_alt_arbiter_acq_2 (
	grant_7,
	mutex_req,
	mutex_grant1)/* synthesis synthesis_greybox=0 */;
input 	grant_7;
input 	mutex_req;
output 	mutex_grant1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb mutex_grant(
	.dataa(!grant_7),
	.datab(!mutex_req),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mutex_grant1),
	.sumout(),
	.cout(),
	.shareout());
defparam mutex_grant.extended_lut = "off";
defparam mutex_grant.lut_mask = 64'h1111111111111111;
defparam mutex_grant.shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_basic_acq_1 (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	ctrl_addr_1,
	ctrl_addr_2,
	ctrl_addr_0,
	ctrl_addr_4,
	ctrl_addr_5,
	ctrl_addr_6,
	ctrl_addr_7,
	ctrl_addr_8,
	ctrl_addr_9,
	ctrl_addr_10,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write1,
	mutex_req1,
	mutex_grant,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read1,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	reset,
	ph_readdata_0,
	logical_ch_addr,
	ph_readdata_1,
	ph_readdata_2,
	ph_readdata_3,
	ph_readdata_4,
	ph_readdata_5,
	ph_readdata_6,
	ph_readdata_7,
	ph_readdata_8,
	ph_readdata_9,
	illegal_phy_ch1,
	ph_readdata_10,
	ph_readdata_11,
	ph_readdata_12,
	ph_readdata_13,
	ph_readdata_14,
	ph_readdata_15,
	ph_readdata_16,
	ph_readdata_17,
	ph_readdata_18,
	ph_readdata_19,
	ph_readdata_20,
	ph_readdata_21,
	ph_readdata_22,
	ph_readdata_23,
	ph_readdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	ctrl_opcode_1,
	ctrl_opcode_2,
	ctrl_opcode_0,
	ctrl_go,
	ctrl_lock,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	waitrequest_to_ctrl1,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	readdata_for_user_0,
	readdata_for_user_1,
	readdata_for_user_2,
	readdata_for_user_3,
	readdata_for_user_4,
	readdata_for_user_5,
	readdata_for_user_6,
	readdata_for_user_7,
	readdata_for_user_8,
	readdata_for_user_9,
	readdata_for_user_10,
	readdata_for_user_11,
	readdata_for_user_12,
	readdata_for_user_13,
	readdata_for_user_14,
	readdata_for_user_15,
	readdata_for_user_16,
	readdata_for_user_17,
	readdata_for_user_18,
	readdata_for_user_19,
	readdata_for_user_20,
	readdata_for_user_21,
	readdata_for_user_22,
	readdata_for_user_23,
	readdata_for_user_24,
	readdata_for_user_25,
	readdata_for_user_26,
	readdata_for_user_27,
	readdata_for_user_28,
	readdata_for_user_29,
	readdata_for_user_30,
	readdata_for_user_31,
	ctrl_wdata_1,
	ctrl_wdata_2,
	ctrl_wdata_0,
	ctrl_wdata_3,
	ctrl_addr_3,
	ctrl_wdata_4,
	ctrl_wdata_5,
	ctrl_wdata_6,
	ctrl_wdata_7,
	ctrl_wdata_8,
	ctrl_wdata_9,
	ctrl_wdata_10,
	ctrl_wdata_11,
	ctrl_addr_11,
	ctrl_wdata_12,
	ctrl_wdata_13,
	ctrl_wdata_14,
	ctrl_wdata_15,
	clk)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_16;
input 	basic_reconfig_readdata_17;
input 	basic_reconfig_readdata_18;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
input 	ctrl_addr_1;
input 	ctrl_addr_2;
input 	ctrl_addr_0;
input 	ctrl_addr_4;
input 	ctrl_addr_5;
input 	ctrl_addr_6;
input 	ctrl_addr_7;
input 	ctrl_addr_8;
input 	ctrl_addr_9;
input 	ctrl_addr_10;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write1;
output 	mutex_req1;
input 	mutex_grant;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read1;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	reset;
output 	ph_readdata_0;
input 	[9:0] logical_ch_addr;
output 	ph_readdata_1;
output 	ph_readdata_2;
output 	ph_readdata_3;
output 	ph_readdata_4;
output 	ph_readdata_5;
output 	ph_readdata_6;
output 	ph_readdata_7;
output 	ph_readdata_8;
output 	ph_readdata_9;
output 	illegal_phy_ch1;
output 	ph_readdata_10;
output 	ph_readdata_11;
output 	ph_readdata_12;
output 	ph_readdata_13;
output 	ph_readdata_14;
output 	ph_readdata_15;
output 	ph_readdata_16;
output 	ph_readdata_17;
output 	ph_readdata_18;
output 	ph_readdata_19;
output 	ph_readdata_20;
output 	ph_readdata_21;
output 	ph_readdata_22;
output 	ph_readdata_23;
output 	ph_readdata_24;
output 	ph_readdata_25;
output 	ph_readdata_26;
output 	ph_readdata_27;
output 	ph_readdata_28;
output 	ph_readdata_29;
output 	ph_readdata_30;
output 	ph_readdata_31;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
input 	ctrl_opcode_1;
input 	ctrl_opcode_2;
input 	ctrl_opcode_0;
input 	ctrl_go;
input 	ctrl_lock;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	waitrequest_to_ctrl1;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
output 	readdata_for_user_0;
output 	readdata_for_user_1;
output 	readdata_for_user_2;
output 	readdata_for_user_3;
output 	readdata_for_user_4;
output 	readdata_for_user_5;
output 	readdata_for_user_6;
output 	readdata_for_user_7;
output 	readdata_for_user_8;
output 	readdata_for_user_9;
output 	readdata_for_user_10;
output 	readdata_for_user_11;
output 	readdata_for_user_12;
output 	readdata_for_user_13;
output 	readdata_for_user_14;
output 	readdata_for_user_15;
output 	readdata_for_user_16;
output 	readdata_for_user_17;
output 	readdata_for_user_18;
output 	readdata_for_user_19;
output 	readdata_for_user_20;
output 	readdata_for_user_21;
output 	readdata_for_user_22;
output 	readdata_for_user_23;
output 	readdata_for_user_24;
output 	readdata_for_user_25;
output 	readdata_for_user_26;
output 	readdata_for_user_27;
output 	readdata_for_user_28;
output 	readdata_for_user_29;
output 	readdata_for_user_30;
output 	readdata_for_user_31;
input 	ctrl_wdata_1;
input 	ctrl_wdata_2;
input 	ctrl_wdata_0;
input 	ctrl_wdata_3;
input 	ctrl_addr_3;
input 	ctrl_wdata_4;
input 	ctrl_wdata_5;
input 	ctrl_wdata_6;
input 	ctrl_wdata_7;
input 	ctrl_wdata_8;
input 	ctrl_wdata_9;
input 	ctrl_wdata_10;
input 	ctrl_wdata_11;
input 	ctrl_addr_11;
input 	ctrl_wdata_12;
input 	ctrl_wdata_13;
input 	ctrl_wdata_14;
input 	ctrl_wdata_15;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state.ST_READ_RECONFIG_BASIC_DATA~q ;
wire \Selector3~3_combout ;
wire \lch_dly[9]~q ;
wire \lch_dly[7]~q ;
wire \lch_dly[8]~q ;
wire \lch_legal~0_combout ;
wire \lch_dly[6]~q ;
wire \lch_dly[4]~q ;
wire \lch_dly[5]~q ;
wire \lch_legal~1_combout ;
wire \Equal2~0_combout ;
wire \lch_dly[0]~q ;
wire \lch_dly[3]~q ;
wire \lch_dly[1]~q ;
wire \lch_dly[2]~q ;
wire \lch_legal~2_combout ;
wire \lch_legal~3_combout ;
wire \lch_legal~4_combout ;
wire \lch_legal~5_combout ;
wire \lch_legal~6_combout ;
wire \lch_legal~q ;
wire \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ;
wire \Selector13~0_combout ;
wire \state.ST_START_AGAIN~q ;
wire \WideOr2~combout ;
wire \Selector3~11_combout ;
wire \Selector3~16_combout ;
wire \Selector3~13_combout ;
wire \Selector15~0_combout ;
wire \Selector10~0_combout ;
wire \Selector15~2_combout ;
wire \phy_addr_is_set~0_combout ;
wire \phy_addr_is_set~q ;
wire \Selector3~8_combout ;
wire \Selector3~9_combout ;
wire \Selector3~10_combout ;
wire \Selector3~12_combout ;
wire \Selector8~0_combout ;
wire \Selector3~17_combout ;
wire \Selector8~1_combout ;
wire \state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ;
wire \Selector9~0_combout ;
wire \state.ST_SET_RECONFIG_BASIC_WRITE~q ;
wire \Selector12~0_combout ;
wire \Selector12~1_combout ;
wire \Selector12~2_combout ;
wire \state.ST_CHECK_CTRLLOCK~q ;
wire \Selector14~0_combout ;
wire \Selector14~1_combout ;
wire \state.ST_RELEASE_REQ~q ;
wire \Selector1~0_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \state.0000~q ;
wire \Selector1~1_combout ;
wire \state.ST_REQ_MUTEX~q ;
wire \Selector2~0_combout ;
wire \state.ST_WRITE_RECONFIG_BASIC_LCH~q ;
wire \Selector3~4_combout ;
wire \Selector3~6_combout ;
wire \state.ST_READ_PHY_ADDRESS~q ;
wire \Selector4~0_combout ;
wire \state.ST_CHECK_PHY_ADD_LEGAL~q ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ;
wire \Selector3~5_combout ;
wire \Selector3~15_combout ;
wire \Selector5~0_combout ;
wire \state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ;
wire \Selector3~7_combout ;
wire \Selector3~14_combout ;
wire \Selector10~1_combout ;
wire \state.ST_SET_RECONFIG_BASIC_READ~q ;
wire \Selector11~0_combout ;
wire \WideOr7~0_combout ;
wire \WideOr8~combout ;
wire \Selector15~1_combout ;
wire \WideOr6~0_combout ;
wire \WideOr5~0_combout ;
wire \WideOr5~1_combout ;
wire \WideOr17~0_combout ;
wire \Selector29~0_combout ;
wire \WideOr7~combout ;
wire \WideOr6~combout ;
wire \WideOr9~combout ;
wire \WideOr17~1_combout ;
wire \WideOr17~2_combout ;
wire \Selector16~0_combout ;
wire \Selector12~3_combout ;
wire \ph_readdata[13]~0_combout ;
wire \ph_readdata[13]~1_combout ;
wire \Selector27~0_combout ;
wire \Selector27~1_combout ;
wire \Selector27~2_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \Selector28~0_combout ;
wire \Selector28~1_combout ;
wire \Selector25~0_combout ;
wire \Selector25~1_combout ;
wire \Selector25~2_combout ;
wire \Selector16~1_combout ;
wire \master_writedata[5]~0_combout ;
wire \master_writedata[5]~1_combout ;
wire \master_writedata[5]~2_combout ;
wire \Selector24~0_combout ;
wire \Selector23~0_combout ;
wire \Selector22~0_combout ;
wire \Selector21~0_combout ;
wire \Selector20~0_combout ;
wire \Selector19~0_combout ;
wire \Selector18~0_combout ;
wire \Selector17~0_combout ;
wire \master_writedata~3_combout ;
wire \master_writedata~4_combout ;
wire \master_writedata~5_combout ;
wire \master_writedata~6_combout ;
wire \readdata_for_user[0]~0_combout ;


dffeas master_write(
	.clk(clk),
	.d(\WideOr8~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write1),
	.prn(vcc));
defparam master_write.is_wysiwyg = "true";
defparam master_write.power_up = "low";

dffeas mutex_req(
	.clk(clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mutex_req1),
	.prn(vcc));
defparam mutex_req.is_wysiwyg = "true";
defparam mutex_req.power_up = "low";

dffeas \master_address[2] (
	.clk(clk),
	.d(\WideOr5~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_2),
	.prn(vcc));
defparam \master_address[2] .is_wysiwyg = "true";
defparam \master_address[2] .power_up = "low";

dffeas \master_address[0] (
	.clk(clk),
	.d(\WideOr7~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_0),
	.prn(vcc));
defparam \master_address[0] .is_wysiwyg = "true";
defparam \master_address[0] .power_up = "low";

dffeas \master_address[1] (
	.clk(clk),
	.d(\WideOr6~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_1),
	.prn(vcc));
defparam \master_address[1] .is_wysiwyg = "true";
defparam \master_address[1] .power_up = "low";

dffeas master_read(
	.clk(clk),
	.d(\WideOr9~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_read1),
	.prn(vcc));
defparam master_read.is_wysiwyg = "true";
defparam master_read.power_up = "low";

dffeas \ph_readdata[0] (
	.clk(clk),
	.d(basic_reconfig_readdata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_0),
	.prn(vcc));
defparam \ph_readdata[0] .is_wysiwyg = "true";
defparam \ph_readdata[0] .power_up = "low";

dffeas \ph_readdata[1] (
	.clk(clk),
	.d(basic_reconfig_readdata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_1),
	.prn(vcc));
defparam \ph_readdata[1] .is_wysiwyg = "true";
defparam \ph_readdata[1] .power_up = "low";

dffeas \ph_readdata[2] (
	.clk(clk),
	.d(basic_reconfig_readdata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_2),
	.prn(vcc));
defparam \ph_readdata[2] .is_wysiwyg = "true";
defparam \ph_readdata[2] .power_up = "low";

dffeas \ph_readdata[3] (
	.clk(clk),
	.d(basic_reconfig_readdata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_3),
	.prn(vcc));
defparam \ph_readdata[3] .is_wysiwyg = "true";
defparam \ph_readdata[3] .power_up = "low";

dffeas \ph_readdata[4] (
	.clk(clk),
	.d(basic_reconfig_readdata_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_4),
	.prn(vcc));
defparam \ph_readdata[4] .is_wysiwyg = "true";
defparam \ph_readdata[4] .power_up = "low";

dffeas \ph_readdata[5] (
	.clk(clk),
	.d(basic_reconfig_readdata_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_5),
	.prn(vcc));
defparam \ph_readdata[5] .is_wysiwyg = "true";
defparam \ph_readdata[5] .power_up = "low";

dffeas \ph_readdata[6] (
	.clk(clk),
	.d(basic_reconfig_readdata_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_6),
	.prn(vcc));
defparam \ph_readdata[6] .is_wysiwyg = "true";
defparam \ph_readdata[6] .power_up = "low";

dffeas \ph_readdata[7] (
	.clk(clk),
	.d(basic_reconfig_readdata_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_7),
	.prn(vcc));
defparam \ph_readdata[7] .is_wysiwyg = "true";
defparam \ph_readdata[7] .power_up = "low";

dffeas \ph_readdata[8] (
	.clk(clk),
	.d(basic_reconfig_readdata_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_8),
	.prn(vcc));
defparam \ph_readdata[8] .is_wysiwyg = "true";
defparam \ph_readdata[8] .power_up = "low";

dffeas \ph_readdata[9] (
	.clk(clk),
	.d(basic_reconfig_readdata_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_9),
	.prn(vcc));
defparam \ph_readdata[9] .is_wysiwyg = "true";
defparam \ph_readdata[9] .power_up = "low";

dffeas illegal_phy_ch(
	.clk(clk),
	.d(Equal8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(illegal_phy_ch1),
	.prn(vcc));
defparam illegal_phy_ch.is_wysiwyg = "true";
defparam illegal_phy_ch.power_up = "low";

dffeas \ph_readdata[10] (
	.clk(clk),
	.d(basic_reconfig_readdata_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_10),
	.prn(vcc));
defparam \ph_readdata[10] .is_wysiwyg = "true";
defparam \ph_readdata[10] .power_up = "low";

dffeas \ph_readdata[11] (
	.clk(clk),
	.d(basic_reconfig_readdata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_11),
	.prn(vcc));
defparam \ph_readdata[11] .is_wysiwyg = "true";
defparam \ph_readdata[11] .power_up = "low";

dffeas \ph_readdata[12] (
	.clk(clk),
	.d(basic_reconfig_readdata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_12),
	.prn(vcc));
defparam \ph_readdata[12] .is_wysiwyg = "true";
defparam \ph_readdata[12] .power_up = "low";

dffeas \ph_readdata[13] (
	.clk(clk),
	.d(basic_reconfig_readdata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_13),
	.prn(vcc));
defparam \ph_readdata[13] .is_wysiwyg = "true";
defparam \ph_readdata[13] .power_up = "low";

dffeas \ph_readdata[14] (
	.clk(clk),
	.d(basic_reconfig_readdata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_14),
	.prn(vcc));
defparam \ph_readdata[14] .is_wysiwyg = "true";
defparam \ph_readdata[14] .power_up = "low";

dffeas \ph_readdata[15] (
	.clk(clk),
	.d(basic_reconfig_readdata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_15),
	.prn(vcc));
defparam \ph_readdata[15] .is_wysiwyg = "true";
defparam \ph_readdata[15] .power_up = "low";

dffeas \ph_readdata[16] (
	.clk(clk),
	.d(basic_reconfig_readdata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_16),
	.prn(vcc));
defparam \ph_readdata[16] .is_wysiwyg = "true";
defparam \ph_readdata[16] .power_up = "low";

dffeas \ph_readdata[17] (
	.clk(clk),
	.d(basic_reconfig_readdata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_17),
	.prn(vcc));
defparam \ph_readdata[17] .is_wysiwyg = "true";
defparam \ph_readdata[17] .power_up = "low";

dffeas \ph_readdata[18] (
	.clk(clk),
	.d(basic_reconfig_readdata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_18),
	.prn(vcc));
defparam \ph_readdata[18] .is_wysiwyg = "true";
defparam \ph_readdata[18] .power_up = "low";

dffeas \ph_readdata[19] (
	.clk(clk),
	.d(basic_reconfig_readdata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_19),
	.prn(vcc));
defparam \ph_readdata[19] .is_wysiwyg = "true";
defparam \ph_readdata[19] .power_up = "low";

dffeas \ph_readdata[20] (
	.clk(clk),
	.d(basic_reconfig_readdata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_20),
	.prn(vcc));
defparam \ph_readdata[20] .is_wysiwyg = "true";
defparam \ph_readdata[20] .power_up = "low";

dffeas \ph_readdata[21] (
	.clk(clk),
	.d(basic_reconfig_readdata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_21),
	.prn(vcc));
defparam \ph_readdata[21] .is_wysiwyg = "true";
defparam \ph_readdata[21] .power_up = "low";

dffeas \ph_readdata[22] (
	.clk(clk),
	.d(basic_reconfig_readdata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_22),
	.prn(vcc));
defparam \ph_readdata[22] .is_wysiwyg = "true";
defparam \ph_readdata[22] .power_up = "low";

dffeas \ph_readdata[23] (
	.clk(clk),
	.d(basic_reconfig_readdata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_23),
	.prn(vcc));
defparam \ph_readdata[23] .is_wysiwyg = "true";
defparam \ph_readdata[23] .power_up = "low";

dffeas \ph_readdata[24] (
	.clk(clk),
	.d(basic_reconfig_readdata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_24),
	.prn(vcc));
defparam \ph_readdata[24] .is_wysiwyg = "true";
defparam \ph_readdata[24] .power_up = "low";

dffeas \ph_readdata[25] (
	.clk(clk),
	.d(basic_reconfig_readdata_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_25),
	.prn(vcc));
defparam \ph_readdata[25] .is_wysiwyg = "true";
defparam \ph_readdata[25] .power_up = "low";

dffeas \ph_readdata[26] (
	.clk(clk),
	.d(basic_reconfig_readdata_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_26),
	.prn(vcc));
defparam \ph_readdata[26] .is_wysiwyg = "true";
defparam \ph_readdata[26] .power_up = "low";

dffeas \ph_readdata[27] (
	.clk(clk),
	.d(basic_reconfig_readdata_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_27),
	.prn(vcc));
defparam \ph_readdata[27] .is_wysiwyg = "true";
defparam \ph_readdata[27] .power_up = "low";

dffeas \ph_readdata[28] (
	.clk(clk),
	.d(basic_reconfig_readdata_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_28),
	.prn(vcc));
defparam \ph_readdata[28] .is_wysiwyg = "true";
defparam \ph_readdata[28] .power_up = "low";

dffeas \ph_readdata[29] (
	.clk(clk),
	.d(basic_reconfig_readdata_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_29),
	.prn(vcc));
defparam \ph_readdata[29] .is_wysiwyg = "true";
defparam \ph_readdata[29] .power_up = "low";

dffeas \ph_readdata[30] (
	.clk(clk),
	.d(basic_reconfig_readdata_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_30),
	.prn(vcc));
defparam \ph_readdata[30] .is_wysiwyg = "true";
defparam \ph_readdata[30] .power_up = "low";

dffeas \ph_readdata[31] (
	.clk(clk),
	.d(basic_reconfig_readdata_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_31),
	.prn(vcc));
defparam \ph_readdata[31] .is_wysiwyg = "true";
defparam \ph_readdata[31] .power_up = "low";

dffeas \master_writedata[1] (
	.clk(clk),
	.d(\Selector27~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_1),
	.prn(vcc));
defparam \master_writedata[1] .is_wysiwyg = "true";
defparam \master_writedata[1] .power_up = "low";

dffeas \master_writedata[2] (
	.clk(clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_2),
	.prn(vcc));
defparam \master_writedata[2] .is_wysiwyg = "true";
defparam \master_writedata[2] .power_up = "low";

dffeas \master_writedata[0] (
	.clk(clk),
	.d(\Selector28~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_0),
	.prn(vcc));
defparam \master_writedata[0] .is_wysiwyg = "true";
defparam \master_writedata[0] .power_up = "low";

dffeas \master_writedata[3] (
	.clk(clk),
	.d(\Selector25~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_3),
	.prn(vcc));
defparam \master_writedata[3] .is_wysiwyg = "true";
defparam \master_writedata[3] .power_up = "low";

dffeas waitrequest_to_ctrl(
	.clk(clk),
	.d(\Selector16~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_to_ctrl1),
	.prn(vcc));
defparam waitrequest_to_ctrl.is_wysiwyg = "true";
defparam waitrequest_to_ctrl.power_up = "low";

dffeas \master_writedata[4] (
	.clk(clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_4),
	.prn(vcc));
defparam \master_writedata[4] .is_wysiwyg = "true";
defparam \master_writedata[4] .power_up = "low";

dffeas \master_writedata[5] (
	.clk(clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_5),
	.prn(vcc));
defparam \master_writedata[5] .is_wysiwyg = "true";
defparam \master_writedata[5] .power_up = "low";

dffeas \master_writedata[6] (
	.clk(clk),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_6),
	.prn(vcc));
defparam \master_writedata[6] .is_wysiwyg = "true";
defparam \master_writedata[6] .power_up = "low";

dffeas \master_writedata[7] (
	.clk(clk),
	.d(\Selector21~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_7),
	.prn(vcc));
defparam \master_writedata[7] .is_wysiwyg = "true";
defparam \master_writedata[7] .power_up = "low";

dffeas \master_writedata[8] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_8),
	.prn(vcc));
defparam \master_writedata[8] .is_wysiwyg = "true";
defparam \master_writedata[8] .power_up = "low";

dffeas \master_writedata[9] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_9),
	.prn(vcc));
defparam \master_writedata[9] .is_wysiwyg = "true";
defparam \master_writedata[9] .power_up = "low";

dffeas \master_writedata[10] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_10),
	.prn(vcc));
defparam \master_writedata[10] .is_wysiwyg = "true";
defparam \master_writedata[10] .power_up = "low";

dffeas \master_writedata[11] (
	.clk(clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_11),
	.prn(vcc));
defparam \master_writedata[11] .is_wysiwyg = "true";
defparam \master_writedata[11] .power_up = "low";

dffeas \master_writedata[12] (
	.clk(clk),
	.d(\master_writedata~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_12),
	.prn(vcc));
defparam \master_writedata[12] .is_wysiwyg = "true";
defparam \master_writedata[12] .power_up = "low";

dffeas \master_writedata[13] (
	.clk(clk),
	.d(\master_writedata~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_13),
	.prn(vcc));
defparam \master_writedata[13] .is_wysiwyg = "true";
defparam \master_writedata[13] .power_up = "low";

dffeas \master_writedata[14] (
	.clk(clk),
	.d(\master_writedata~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_14),
	.prn(vcc));
defparam \master_writedata[14] .is_wysiwyg = "true";
defparam \master_writedata[14] .power_up = "low";

dffeas \master_writedata[15] (
	.clk(clk),
	.d(\master_writedata~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_15),
	.prn(vcc));
defparam \master_writedata[15] .is_wysiwyg = "true";
defparam \master_writedata[15] .power_up = "low";

dffeas \readdata_for_user[0] (
	.clk(clk),
	.d(basic_reconfig_readdata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_0),
	.prn(vcc));
defparam \readdata_for_user[0] .is_wysiwyg = "true";
defparam \readdata_for_user[0] .power_up = "low";

dffeas \readdata_for_user[1] (
	.clk(clk),
	.d(basic_reconfig_readdata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_1),
	.prn(vcc));
defparam \readdata_for_user[1] .is_wysiwyg = "true";
defparam \readdata_for_user[1] .power_up = "low";

dffeas \readdata_for_user[2] (
	.clk(clk),
	.d(basic_reconfig_readdata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_2),
	.prn(vcc));
defparam \readdata_for_user[2] .is_wysiwyg = "true";
defparam \readdata_for_user[2] .power_up = "low";

dffeas \readdata_for_user[3] (
	.clk(clk),
	.d(basic_reconfig_readdata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_3),
	.prn(vcc));
defparam \readdata_for_user[3] .is_wysiwyg = "true";
defparam \readdata_for_user[3] .power_up = "low";

dffeas \readdata_for_user[4] (
	.clk(clk),
	.d(basic_reconfig_readdata_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_4),
	.prn(vcc));
defparam \readdata_for_user[4] .is_wysiwyg = "true";
defparam \readdata_for_user[4] .power_up = "low";

dffeas \readdata_for_user[5] (
	.clk(clk),
	.d(basic_reconfig_readdata_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_5),
	.prn(vcc));
defparam \readdata_for_user[5] .is_wysiwyg = "true";
defparam \readdata_for_user[5] .power_up = "low";

dffeas \readdata_for_user[6] (
	.clk(clk),
	.d(basic_reconfig_readdata_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_6),
	.prn(vcc));
defparam \readdata_for_user[6] .is_wysiwyg = "true";
defparam \readdata_for_user[6] .power_up = "low";

dffeas \readdata_for_user[7] (
	.clk(clk),
	.d(basic_reconfig_readdata_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_7),
	.prn(vcc));
defparam \readdata_for_user[7] .is_wysiwyg = "true";
defparam \readdata_for_user[7] .power_up = "low";

dffeas \readdata_for_user[8] (
	.clk(clk),
	.d(basic_reconfig_readdata_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_8),
	.prn(vcc));
defparam \readdata_for_user[8] .is_wysiwyg = "true";
defparam \readdata_for_user[8] .power_up = "low";

dffeas \readdata_for_user[9] (
	.clk(clk),
	.d(basic_reconfig_readdata_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_9),
	.prn(vcc));
defparam \readdata_for_user[9] .is_wysiwyg = "true";
defparam \readdata_for_user[9] .power_up = "low";

dffeas \readdata_for_user[10] (
	.clk(clk),
	.d(basic_reconfig_readdata_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_10),
	.prn(vcc));
defparam \readdata_for_user[10] .is_wysiwyg = "true";
defparam \readdata_for_user[10] .power_up = "low";

dffeas \readdata_for_user[11] (
	.clk(clk),
	.d(basic_reconfig_readdata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_11),
	.prn(vcc));
defparam \readdata_for_user[11] .is_wysiwyg = "true";
defparam \readdata_for_user[11] .power_up = "low";

dffeas \readdata_for_user[12] (
	.clk(clk),
	.d(basic_reconfig_readdata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_12),
	.prn(vcc));
defparam \readdata_for_user[12] .is_wysiwyg = "true";
defparam \readdata_for_user[12] .power_up = "low";

dffeas \readdata_for_user[13] (
	.clk(clk),
	.d(basic_reconfig_readdata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_13),
	.prn(vcc));
defparam \readdata_for_user[13] .is_wysiwyg = "true";
defparam \readdata_for_user[13] .power_up = "low";

dffeas \readdata_for_user[14] (
	.clk(clk),
	.d(basic_reconfig_readdata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_14),
	.prn(vcc));
defparam \readdata_for_user[14] .is_wysiwyg = "true";
defparam \readdata_for_user[14] .power_up = "low";

dffeas \readdata_for_user[15] (
	.clk(clk),
	.d(basic_reconfig_readdata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_15),
	.prn(vcc));
defparam \readdata_for_user[15] .is_wysiwyg = "true";
defparam \readdata_for_user[15] .power_up = "low";

dffeas \readdata_for_user[16] (
	.clk(clk),
	.d(basic_reconfig_readdata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_16),
	.prn(vcc));
defparam \readdata_for_user[16] .is_wysiwyg = "true";
defparam \readdata_for_user[16] .power_up = "low";

dffeas \readdata_for_user[17] (
	.clk(clk),
	.d(basic_reconfig_readdata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_17),
	.prn(vcc));
defparam \readdata_for_user[17] .is_wysiwyg = "true";
defparam \readdata_for_user[17] .power_up = "low";

dffeas \readdata_for_user[18] (
	.clk(clk),
	.d(basic_reconfig_readdata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_18),
	.prn(vcc));
defparam \readdata_for_user[18] .is_wysiwyg = "true";
defparam \readdata_for_user[18] .power_up = "low";

dffeas \readdata_for_user[19] (
	.clk(clk),
	.d(basic_reconfig_readdata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_19),
	.prn(vcc));
defparam \readdata_for_user[19] .is_wysiwyg = "true";
defparam \readdata_for_user[19] .power_up = "low";

dffeas \readdata_for_user[20] (
	.clk(clk),
	.d(basic_reconfig_readdata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_20),
	.prn(vcc));
defparam \readdata_for_user[20] .is_wysiwyg = "true";
defparam \readdata_for_user[20] .power_up = "low";

dffeas \readdata_for_user[21] (
	.clk(clk),
	.d(basic_reconfig_readdata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_21),
	.prn(vcc));
defparam \readdata_for_user[21] .is_wysiwyg = "true";
defparam \readdata_for_user[21] .power_up = "low";

dffeas \readdata_for_user[22] (
	.clk(clk),
	.d(basic_reconfig_readdata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_22),
	.prn(vcc));
defparam \readdata_for_user[22] .is_wysiwyg = "true";
defparam \readdata_for_user[22] .power_up = "low";

dffeas \readdata_for_user[23] (
	.clk(clk),
	.d(basic_reconfig_readdata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_23),
	.prn(vcc));
defparam \readdata_for_user[23] .is_wysiwyg = "true";
defparam \readdata_for_user[23] .power_up = "low";

dffeas \readdata_for_user[24] (
	.clk(clk),
	.d(basic_reconfig_readdata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_24),
	.prn(vcc));
defparam \readdata_for_user[24] .is_wysiwyg = "true";
defparam \readdata_for_user[24] .power_up = "low";

dffeas \readdata_for_user[25] (
	.clk(clk),
	.d(basic_reconfig_readdata_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_25),
	.prn(vcc));
defparam \readdata_for_user[25] .is_wysiwyg = "true";
defparam \readdata_for_user[25] .power_up = "low";

dffeas \readdata_for_user[26] (
	.clk(clk),
	.d(basic_reconfig_readdata_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_26),
	.prn(vcc));
defparam \readdata_for_user[26] .is_wysiwyg = "true";
defparam \readdata_for_user[26] .power_up = "low";

dffeas \readdata_for_user[27] (
	.clk(clk),
	.d(basic_reconfig_readdata_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_27),
	.prn(vcc));
defparam \readdata_for_user[27] .is_wysiwyg = "true";
defparam \readdata_for_user[27] .power_up = "low";

dffeas \readdata_for_user[28] (
	.clk(clk),
	.d(basic_reconfig_readdata_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_28),
	.prn(vcc));
defparam \readdata_for_user[28] .is_wysiwyg = "true";
defparam \readdata_for_user[28] .power_up = "low";

dffeas \readdata_for_user[29] (
	.clk(clk),
	.d(basic_reconfig_readdata_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_29),
	.prn(vcc));
defparam \readdata_for_user[29] .is_wysiwyg = "true";
defparam \readdata_for_user[29] .power_up = "low";

dffeas \readdata_for_user[30] (
	.clk(clk),
	.d(basic_reconfig_readdata_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_30),
	.prn(vcc));
defparam \readdata_for_user[30] .is_wysiwyg = "true";
defparam \readdata_for_user[30] .power_up = "low";

dffeas \readdata_for_user[31] (
	.clk(clk),
	.d(basic_reconfig_readdata_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_31),
	.prn(vcc));
defparam \readdata_for_user[31] .is_wysiwyg = "true";
defparam \readdata_for_user[31] .power_up = "low";

dffeas \state.ST_READ_RECONFIG_BASIC_DATA (
	.clk(clk),
	.d(\Selector11~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.prn(vcc));
defparam \state.ST_READ_RECONFIG_BASIC_DATA .is_wysiwyg = "true";
defparam \state.ST_READ_RECONFIG_BASIC_DATA .power_up = "low";

cyclonev_lcell_comb \Selector3~3 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!basic_reconfig_readdata_1),
	.datac(!basic_reconfig_readdata_2),
	.datad(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~3 .extended_lut = "off";
defparam \Selector3~3 .lut_mask = 64'h0001000100010001;
defparam \Selector3~3 .shared_arith = "off";

dffeas \lch_dly[9] (
	.clk(clk),
	.d(logical_ch_addr[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[9]~q ),
	.prn(vcc));
defparam \lch_dly[9] .is_wysiwyg = "true";
defparam \lch_dly[9] .power_up = "low";

dffeas \lch_dly[7] (
	.clk(clk),
	.d(logical_ch_addr[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[7]~q ),
	.prn(vcc));
defparam \lch_dly[7] .is_wysiwyg = "true";
defparam \lch_dly[7] .power_up = "low";

dffeas \lch_dly[8] (
	.clk(clk),
	.d(logical_ch_addr[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[8]~q ),
	.prn(vcc));
defparam \lch_dly[8] .is_wysiwyg = "true";
defparam \lch_dly[8] .power_up = "low";

cyclonev_lcell_comb \lch_legal~0 (
	.dataa(!logical_ch_addr[7]),
	.datab(!logical_ch_addr[8]),
	.datac(!\lch_dly[7]~q ),
	.datad(!\lch_dly[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~0 .extended_lut = "off";
defparam \lch_legal~0 .lut_mask = 64'h8421842184218421;
defparam \lch_legal~0 .shared_arith = "off";

dffeas \lch_dly[6] (
	.clk(clk),
	.d(logical_ch_addr[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[6]~q ),
	.prn(vcc));
defparam \lch_dly[6] .is_wysiwyg = "true";
defparam \lch_dly[6] .power_up = "low";

dffeas \lch_dly[4] (
	.clk(clk),
	.d(logical_ch_addr[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[4]~q ),
	.prn(vcc));
defparam \lch_dly[4] .is_wysiwyg = "true";
defparam \lch_dly[4] .power_up = "low";

dffeas \lch_dly[5] (
	.clk(clk),
	.d(logical_ch_addr[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[5]~q ),
	.prn(vcc));
defparam \lch_dly[5] .is_wysiwyg = "true";
defparam \lch_dly[5] .power_up = "low";

cyclonev_lcell_comb \lch_legal~1 (
	.dataa(!logical_ch_addr[4]),
	.datab(!logical_ch_addr[5]),
	.datac(!\lch_dly[4]~q ),
	.datad(!\lch_dly[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~1 .extended_lut = "off";
defparam \lch_legal~1 .lut_mask = 64'h8421842184218421;
defparam \lch_legal~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_2),
	.datac(!ctrl_opcode_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h4040404040404040;
defparam \Equal2~0 .shared_arith = "off";

dffeas \lch_dly[0] (
	.clk(clk),
	.d(logical_ch_addr[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[0]~q ),
	.prn(vcc));
defparam \lch_dly[0] .is_wysiwyg = "true";
defparam \lch_dly[0] .power_up = "low";

dffeas \lch_dly[3] (
	.clk(clk),
	.d(logical_ch_addr[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[3]~q ),
	.prn(vcc));
defparam \lch_dly[3] .is_wysiwyg = "true";
defparam \lch_dly[3] .power_up = "low";

dffeas \lch_dly[1] (
	.clk(clk),
	.d(logical_ch_addr[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[1]~q ),
	.prn(vcc));
defparam \lch_dly[1] .is_wysiwyg = "true";
defparam \lch_dly[1] .power_up = "low";

dffeas \lch_dly[2] (
	.clk(clk),
	.d(logical_ch_addr[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[2]~q ),
	.prn(vcc));
defparam \lch_dly[2] .is_wysiwyg = "true";
defparam \lch_dly[2] .power_up = "low";

cyclonev_lcell_comb \lch_legal~2 (
	.dataa(!logical_ch_addr[1]),
	.datab(!logical_ch_addr[2]),
	.datac(!\lch_dly[1]~q ),
	.datad(!\lch_dly[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~2 .extended_lut = "off";
defparam \lch_legal~2 .lut_mask = 64'h8421842184218421;
defparam \lch_legal~2 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~3 (
	.dataa(!logical_ch_addr[0]),
	.datab(!logical_ch_addr[3]),
	.datac(!\Equal2~0_combout ),
	.datad(!\lch_dly[0]~q ),
	.datae(!\lch_dly[3]~q ),
	.dataf(!\lch_legal~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~3 .extended_lut = "off";
defparam \lch_legal~3 .lut_mask = 64'h0000000080402010;
defparam \lch_legal~3 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~4 (
	.dataa(!logical_ch_addr[6]),
	.datab(!\lch_dly[6]~q ),
	.datac(!\lch_legal~1_combout ),
	.datad(!\lch_legal~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~4 .extended_lut = "off";
defparam \lch_legal~4 .lut_mask = 64'h0009000900090009;
defparam \lch_legal~4 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~5 (
	.dataa(!logical_ch_addr[9]),
	.datab(!\lch_dly[9]~q ),
	.datac(!\lch_legal~0_combout ),
	.datad(!\lch_legal~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~5 .extended_lut = "off";
defparam \lch_legal~5 .lut_mask = 64'h0009000900090009;
defparam \lch_legal~5 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~6 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!Equal8),
	.datac(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datad(!\lch_legal~q ),
	.datae(!\lch_legal~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~6 .extended_lut = "off";
defparam \lch_legal~6 .lut_mask = 64'h000008FF000008FF;
defparam \lch_legal~6 .shared_arith = "off";

dffeas lch_legal(
	.clk(clk),
	.d(\lch_legal~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_legal~q ),
	.prn(vcc));
defparam lch_legal.is_wysiwyg = "true";
defparam lch_legal.power_up = "low";

dffeas \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE (
	.clk(clk),
	.d(\Selector15~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.prn(vcc));
defparam \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE .is_wysiwyg = "true";
defparam \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE .power_up = "low";

cyclonev_lcell_comb \Selector13~0 (
	.dataa(!ctrl_go),
	.datab(!\state.ST_START_AGAIN~q ),
	.datac(!ctrl_lock),
	.datad(!\state.ST_CHECK_CTRLLOCK~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~0 .extended_lut = "off";
defparam \Selector13~0 .lut_mask = 64'h222F222F222F222F;
defparam \Selector13~0 .shared_arith = "off";

dffeas \state.ST_START_AGAIN (
	.clk(clk),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_START_AGAIN~q ),
	.prn(vcc));
defparam \state.ST_START_AGAIN .is_wysiwyg = "true";
defparam \state.ST_START_AGAIN .power_up = "low";

cyclonev_lcell_comb WideOr2(
	.dataa(!\state.ST_REQ_MUTEX~q ),
	.datab(!\state.0000~q ),
	.datac(!\state.ST_START_AGAIN~q ),
	.datad(!\state.ST_CHECK_CTRLLOCK~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr2~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr2.extended_lut = "off";
defparam WideOr2.lut_mask = 64'h2000200020002000;
defparam WideOr2.shared_arith = "off";

cyclonev_lcell_comb \Selector3~11 (
	.dataa(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datab(!\Selector3~4_combout ),
	.datac(!\Selector3~8_combout ),
	.datad(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~11 .extended_lut = "off";
defparam \Selector3~11 .lut_mask = 64'h8000800080008000;
defparam \Selector3~11 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~16 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\Selector3~3_combout ),
	.datad(!\Selector3~4_combout ),
	.datae(!\WideOr2~combout ),
	.dataf(!\Selector3~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~16 .extended_lut = "off";
defparam \Selector3~16 .lut_mask = 64'h0000000000002000;
defparam \Selector3~16 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~13 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_2),
	.datac(!ctrl_opcode_0),
	.datad(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datae(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~13 .extended_lut = "off";
defparam \Selector3~13 .lut_mask = 64'h00AC121200AC1212;
defparam \Selector3~13 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\WideOr2~combout ),
	.dataf(!\Selector3~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "off";
defparam \Selector15~0 .lut_mask = 64'h0000FFFF00007FFF;
defparam \Selector15~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\Selector3~3_combout ),
	.datad(!\Selector3~4_combout ),
	.datae(!\Selector3~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'hF0D0D0D0F0D0D0D0;
defparam \Selector10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~2 (
	.dataa(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datab(!\Selector3~9_combout ),
	.datac(!\Selector3~16_combout ),
	.datad(!\Selector15~0_combout ),
	.datae(!\Selector10~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~2 .extended_lut = "off";
defparam \Selector15~2 .lut_mask = 64'h0000337300003373;
defparam \Selector15~2 .shared_arith = "off";

cyclonev_lcell_comb \phy_addr_is_set~0 (
	.dataa(!\phy_addr_is_set~q ),
	.datab(!\Selector15~2_combout ),
	.datac(!\Selector5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\phy_addr_is_set~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \phy_addr_is_set~0 .extended_lut = "off";
defparam \phy_addr_is_set~0 .lut_mask = 64'h4C4C4C4C4C4C4C4C;
defparam \phy_addr_is_set~0 .shared_arith = "off";

dffeas phy_addr_is_set(
	.clk(clk),
	.d(\phy_addr_is_set~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\phy_addr_is_set~q ),
	.prn(vcc));
defparam phy_addr_is_set.is_wysiwyg = "true";
defparam phy_addr_is_set.power_up = "low";

cyclonev_lcell_comb \Selector3~8 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.datab(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.datac(!\phy_addr_is_set~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~8 .extended_lut = "off";
defparam \Selector3~8 .lut_mask = 64'h0707070707070707;
defparam \Selector3~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~9 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~9 .extended_lut = "off";
defparam \Selector3~9 .lut_mask = 64'h0000800000008000;
defparam \Selector3~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~10 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~3_combout ),
	.dataf(!\Selector3~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~10 .extended_lut = "off";
defparam \Selector3~10 .lut_mask = 64'hFFFF00007FFF0000;
defparam \Selector3~10 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~12 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~12 .extended_lut = "off";
defparam \Selector3~12 .lut_mask = 64'h0000800000008000;
defparam \Selector3~12 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!\Selector3~15_combout ),
	.datab(!\Selector3~9_combout ),
	.datac(!\Selector3~10_combout ),
	.datad(!\WideOr2~combout ),
	.datae(!\Selector3~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h0008000000080000;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~17 (
	.dataa(!\Selector3~15_combout ),
	.datab(!\Selector3~9_combout ),
	.datac(!\Selector3~10_combout ),
	.datad(!\WideOr2~combout ),
	.datae(!\Selector3~12_combout ),
	.dataf(!\Selector15~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~17 .extended_lut = "off";
defparam \Selector3~17 .lut_mask = 64'h0000000008080800;
defparam \Selector3~17 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~1 (
	.dataa(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datab(!\Selector3~7_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!\Selector3~17_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~1 .extended_lut = "off";
defparam \Selector8~1 .lut_mask = 64'h0355035503550355;
defparam \Selector8~1 .shared_arith = "off";

dffeas \state.ST_WRITE_DATA_TO_RECONFIG_BASIC (
	.clk(clk),
	.d(\Selector8~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.prn(vcc));
defparam \state.ST_WRITE_DATA_TO_RECONFIG_BASIC .is_wysiwyg = "true";
defparam \state.ST_WRITE_DATA_TO_RECONFIG_BASIC .power_up = "low";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.dataf(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h00007FFF8000FFFF;
defparam \Selector9~0 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_WRITE (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_WRITE .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_WRITE .power_up = "low";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.datab(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'h8888888888888888;
defparam \Selector12~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~1 (
	.dataa(!Equal8),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datad(!\Equal2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~1 .extended_lut = "off";
defparam \Selector12~1 .lut_mask = 64'hF0D0F0D0F0D0F0D0;
defparam \Selector12~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~2 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_CHECK_CTRLLOCK~q ),
	.datad(!\Selector12~0_combout ),
	.datae(!\phy_addr_is_set~q ),
	.dataf(!\Selector12~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~2 .extended_lut = "off";
defparam \Selector12~2 .lut_mask = 64'h2F222F222F000D00;
defparam \Selector12~2 .shared_arith = "off";

dffeas \state.ST_CHECK_CTRLLOCK (
	.clk(clk),
	.d(\Selector12~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CHECK_CTRLLOCK~q ),
	.prn(vcc));
defparam \state.ST_CHECK_CTRLLOCK .is_wysiwyg = "true";
defparam \state.ST_CHECK_CTRLLOCK .power_up = "low";

cyclonev_lcell_comb \Selector14~0 (
	.dataa(!ctrl_lock),
	.datab(!\state.ST_CHECK_CTRLLOCK~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~0 .extended_lut = "off";
defparam \Selector14~0 .lut_mask = 64'h2222222222222222;
defparam \Selector14~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector14~1 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_RELEASE_REQ~q ),
	.dataf(!\Selector14~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~1 .extended_lut = "off";
defparam \Selector14~1 .lut_mask = 64'h00007FFFFFFFFFFF;
defparam \Selector14~1 .shared_arith = "off";

dffeas \state.ST_RELEASE_REQ (
	.clk(clk),
	.d(\Selector14~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_RELEASE_REQ~q ),
	.prn(vcc));
defparam \state.ST_RELEASE_REQ .is_wysiwyg = "true";
defparam \state.ST_RELEASE_REQ .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!ctrl_go),
	.datab(!ctrl_opcode_1),
	.datac(!ctrl_opcode_2),
	.datad(!ctrl_opcode_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5554555455545554;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\state.0000~q ),
	.datab(!\Selector1~0_combout ),
	.datac(!\Selector3~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h7070707070707070;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~1 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_RELEASE_REQ~q ),
	.dataf(!\Selector0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~1 .extended_lut = "off";
defparam \Selector0~1 .lut_mask = 64'h00000000FFFF7FFF;
defparam \Selector0~1 .shared_arith = "off";

dffeas \state.0000 (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.0000~q ),
	.prn(vcc));
defparam \state.0000 .is_wysiwyg = "true";
defparam \state.0000 .power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!mutex_grant),
	.datab(!\state.ST_REQ_MUTEX~q ),
	.datac(!\state.0000~q ),
	.datad(!\Selector1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h22F222F222F222F2;
defparam \Selector1~1 .shared_arith = "off";

dffeas \state.ST_REQ_MUTEX (
	.clk(clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_REQ_MUTEX~q ),
	.prn(vcc));
defparam \state.ST_REQ_MUTEX .is_wysiwyg = "true";
defparam \state.ST_REQ_MUTEX .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.ST_REQ_MUTEX~q ),
	.datae(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h0055F3F70055F3F7;
defparam \Selector2~0 .shared_arith = "off";

dffeas \state.ST_WRITE_RECONFIG_BASIC_LCH (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.prn(vcc));
defparam \state.ST_WRITE_RECONFIG_BASIC_LCH .is_wysiwyg = "true";
defparam \state.ST_WRITE_RECONFIG_BASIC_LCH .power_up = "low";

cyclonev_lcell_comb \Selector3~4 (
	.dataa(!\lch_legal~q ),
	.datab(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~4 .extended_lut = "off";
defparam \Selector3~4 .lut_mask = 64'h2222222222222222;
defparam \Selector3~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~6 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\Selector3~3_combout ),
	.datad(!\Selector3~4_combout ),
	.datae(!\state.ST_READ_PHY_ADDRESS~q ),
	.dataf(!\Selector3~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~6 .extended_lut = "off";
defparam \Selector3~6 .lut_mask = 64'h0020D0F00000D0D0;
defparam \Selector3~6 .shared_arith = "off";

dffeas \state.ST_READ_PHY_ADDRESS (
	.clk(clk),
	.d(\Selector3~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_READ_PHY_ADDRESS~q ),
	.prn(vcc));
defparam \state.ST_READ_PHY_ADDRESS .is_wysiwyg = "true";
defparam \state.ST_READ_PHY_ADDRESS .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!Equal8),
	.datac(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datad(!\state.ST_READ_PHY_ADDRESS~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h04AE04AE04AE04AE;
defparam \Selector4~0 .shared_arith = "off";

dffeas \state.ST_CHECK_PHY_ADD_LEGAL (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.prn(vcc));
defparam \state.ST_CHECK_PHY_ADD_LEGAL .is_wysiwyg = "true";
defparam \state.ST_CHECK_PHY_ADD_LEGAL .power_up = "low";

cyclonev_lcell_comb \Selector6~1 (
	.dataa(!Equal8),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!\lch_legal~q ),
	.datad(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datae(!\Equal2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'h222F000F222F000F;
defparam \Selector6~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~2 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.datae(!\Selector6~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~2 .extended_lut = "off";
defparam \Selector6~2 .lut_mask = 64'h00FB0CFF00FB0CFF;
defparam \Selector6~2 .shared_arith = "off";

dffeas \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK (
	.clk(clk),
	.d(\Selector6~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.prn(vcc));
defparam \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK .is_wysiwyg = "true";
defparam \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK .power_up = "low";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!ctrl_go),
	.datab(!ctrl_opcode_1),
	.datac(!ctrl_opcode_2),
	.datad(!ctrl_opcode_0),
	.datae(!\state.ST_START_AGAIN~q ),
	.dataf(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h0000555530037557;
defparam \Selector7~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~1 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datae(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.dataf(!\Selector7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~1 .extended_lut = "off";
defparam \Selector7~1 .lut_mask = 64'h00F304F7FFFFFFFF;
defparam \Selector7~1 .shared_arith = "off";

dffeas \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG (
	.clk(clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.prn(vcc));
defparam \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG .is_wysiwyg = "true";
defparam \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG .power_up = "low";

cyclonev_lcell_comb \Selector3~5 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_2),
	.datac(!ctrl_opcode_0),
	.datad(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~5 .extended_lut = "off";
defparam \Selector3~5 .lut_mask = 64'h0012001200120012;
defparam \Selector3~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~15 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~15 .extended_lut = "off";
defparam \Selector3~15 .lut_mask = 64'h0000800000008000;
defparam \Selector3~15 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!\Selector3~15_combout ),
	.datab(!\Selector3~9_combout ),
	.datac(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.datad(!\Selector3~10_combout ),
	.datae(!\Selector3~16_combout ),
	.dataf(!\Selector15~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h55555555555D5555;
defparam \Selector5~0 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_PADDR_MODE (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_PADDR_MODE .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_PADDR_MODE .power_up = "low";

cyclonev_lcell_comb \Selector3~7 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_2),
	.datac(!ctrl_opcode_0),
	.datad(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~7 .extended_lut = "off";
defparam \Selector3~7 .lut_mask = 64'h0C100C100C100C10;
defparam \Selector3~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~14 (
	.dataa(!\Selector3~9_combout ),
	.datab(!\Selector3~10_combout ),
	.datac(!\WideOr2~combout ),
	.datad(!\Selector3~12_combout ),
	.datae(!\Selector15~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~14 .extended_lut = "off";
defparam \Selector3~14 .lut_mask = 64'h0000AAA80000AAA8;
defparam \Selector3~14 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~1 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.datab(!\Selector3~7_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Selector3~14_combout ),
	.datae(!\Selector8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~1 .extended_lut = "off";
defparam \Selector10~1 .lut_mask = 64'h0005CC050005CC05;
defparam \Selector10~1 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_READ (
	.clk(clk),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_READ .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_READ .power_up = "low";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.dataf(!\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h00007FFF8000FFFF;
defparam \Selector11~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr7~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\Selector13~0_combout ),
	.datac(!\Selector4~0_combout ),
	.datad(!\Selector12~2_combout ),
	.datae(!\Selector3~6_combout ),
	.dataf(!\Selector0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr7~0 .extended_lut = "off";
defparam \WideOr7~0 .lut_mask = 64'h0000000080000000;
defparam \WideOr7~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr8(
	.dataa(!\Selector11~0_combout ),
	.datab(!\Selector6~2_combout ),
	.datac(!\WideOr7~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr8~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr8.extended_lut = "off";
defparam WideOr8.lut_mask = 64'h0808080808080808;
defparam WideOr8.shared_arith = "off";

cyclonev_lcell_comb \Selector15~1 (
	.dataa(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datab(!\Selector3~10_combout ),
	.datac(!\WideOr2~combout ),
	.datad(!\Selector3~12_combout ),
	.datae(!\Selector15~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~1 .extended_lut = "off";
defparam \Selector15~1 .lut_mask = 64'h0000555400005554;
defparam \Selector15~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr6~0 (
	.dataa(!\Selector6~2_combout ),
	.datab(!\Selector3~6_combout ),
	.datac(!\Selector9~0_combout ),
	.datad(!\Selector3~9_combout ),
	.datae(!\Selector15~1_combout ),
	.dataf(!\Selector10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr6~0 .extended_lut = "off";
defparam \WideOr6~0 .lut_mask = 64'h8080808080000000;
defparam \WideOr6~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr5~0 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!basic_reconfig_waitrequest2),
	.datac(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datad(!\Selector11~0_combout ),
	.datae(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.dataf(!\Selector7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr5~0 .extended_lut = "off";
defparam \WideOr5~0 .lut_mask = 64'hFC00B80000000000;
defparam \WideOr5~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr5~1 (
	.dataa(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datab(!\Selector3~7_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!\Selector3~17_combout ),
	.datae(!\WideOr5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr5~1 .extended_lut = "off";
defparam \WideOr5~1 .lut_mask = 64'hFFFF0355FFFF0355;
defparam \WideOr5~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr17~0 (
	.dataa(!\Selector13~0_combout ),
	.datab(!\Selector2~0_combout ),
	.datac(!\Selector10~1_combout ),
	.datad(!\Selector5~0_combout ),
	.datae(!\WideOr6~0_combout ),
	.dataf(!\WideOr5~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~0 .extended_lut = "off";
defparam \WideOr17~0 .lut_mask = 64'h0000800000000000;
defparam \WideOr17~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!mutex_req1),
	.datab(!\Selector1~1_combout ),
	.datac(!\Selector4~0_combout ),
	.datad(!\Selector12~2_combout ),
	.datae(!\WideOr17~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'h7777377777773777;
defparam \Selector29~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr7(
	.dataa(!\WideOr7~0_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr7~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr7.extended_lut = "off";
defparam WideOr7.lut_mask = 64'h4444444444444444;
defparam WideOr7.shared_arith = "off";

cyclonev_lcell_comb WideOr6(
	.dataa(!\Selector10~1_combout ),
	.datab(!\Selector5~0_combout ),
	.datac(!\WideOr6~0_combout ),
	.datad(!\Selector14~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr6~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr6.extended_lut = "off";
defparam WideOr6.lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam WideOr6.shared_arith = "off";

cyclonev_lcell_comb WideOr9(
	.dataa(!\Selector11~0_combout ),
	.datab(!\Selector6~2_combout ),
	.datac(!\Selector3~6_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr9~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr9.extended_lut = "off";
defparam WideOr9.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam WideOr9.shared_arith = "off";

cyclonev_lcell_comb \WideOr17~1 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.ST_REQ_MUTEX~q ),
	.datae(!\Selector13~0_combout ),
	.dataf(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~1 .extended_lut = "off";
defparam \WideOr17~1 .lut_mask = 64'hFFAA00000C080000;
defparam \WideOr17~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr17~2 (
	.dataa(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datab(!\Selector3~7_combout ),
	.datac(!\Selector8~0_combout ),
	.datad(!\Selector3~17_combout ),
	.datae(!\WideOr5~0_combout ),
	.dataf(!\WideOr17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~2 .extended_lut = "off";
defparam \WideOr17~2 .lut_mask = 64'h000000000000FCAA;
defparam \WideOr17~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\Selector1~1_combout ),
	.datad(!\state.ST_RELEASE_REQ~q ),
	.datae(!\Selector14~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'hF0200000F0200000;
defparam \Selector16~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~3 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_CHECK_CTRLLOCK~q ),
	.dataf(!\phy_addr_is_set~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~3 .extended_lut = "off";
defparam \Selector12~3 .lut_mask = 64'h8000FFFF00007FFF;
defparam \Selector12~3 .shared_arith = "off";

cyclonev_lcell_comb \ph_readdata[13]~0 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!\Selector12~0_combout ),
	.datad(!\Selector12~3_combout ),
	.datae(!\Selector12~1_combout ),
	.dataf(!\Selector0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ph_readdata[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ph_readdata[13]~0 .extended_lut = "off";
defparam \ph_readdata[13]~0 .lut_mask = 64'h000000007737FF3F;
defparam \ph_readdata[13]~0 .shared_arith = "off";

cyclonev_lcell_comb \ph_readdata[13]~1 (
	.dataa(!\Selector10~1_combout ),
	.datab(!\Selector5~0_combout ),
	.datac(!\WideOr6~0_combout ),
	.datad(!\WideOr17~2_combout ),
	.datae(!\Selector16~0_combout ),
	.dataf(!\ph_readdata[13]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ph_readdata[13]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ph_readdata[13]~1 .extended_lut = "off";
defparam \ph_readdata[13]~1 .lut_mask = 64'h0000000000000008;
defparam \ph_readdata[13]~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_2),
	.datac(!ctrl_opcode_0),
	.datad(!\Selector10~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h0020002000200020;
defparam \Selector27~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~1 (
	.dataa(!logical_ch_addr[1]),
	.datab(!\Selector2~0_combout ),
	.datac(!\Selector7~1_combout ),
	.datad(!ctrl_addr_1),
	.datae(!\Selector27~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~1 .extended_lut = "off";
defparam \Selector27~1 .lut_mask = 64'hEEE00000EEE00000;
defparam \Selector27~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~2 (
	.dataa(!\Selector15~2_combout ),
	.datab(!\Selector5~0_combout ),
	.datac(!\Selector8~1_combout ),
	.datad(!ctrl_wdata_1),
	.datae(!\Selector27~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~2 .extended_lut = "off";
defparam \Selector27~2 .lut_mask = 64'hFFFF777FFFFF777F;
defparam \Selector27~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!logical_ch_addr[2]),
	.datab(!\Selector2~0_combout ),
	.datac(!\Selector14~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \Selector26~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~1 (
	.dataa(!\Selector8~1_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(!ctrl_wdata_2),
	.datad(!ctrl_addr_2),
	.datae(!\Selector26~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~1 .extended_lut = "off";
defparam \Selector26~1 .lut_mask = 64'hFFFF0537FFFF0537;
defparam \Selector26~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!logical_ch_addr[0]),
	.datab(!\Selector2~0_combout ),
	.datac(!\Selector7~1_combout ),
	.datad(!ctrl_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h111F111F111F111F;
defparam \Selector28~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~1 (
	.dataa(!\Selector10~1_combout ),
	.datab(!\Selector5~0_combout ),
	.datac(!\Selector8~1_combout ),
	.datad(!ctrl_wdata_0),
	.datae(!\Selector28~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~1 .extended_lut = "off";
defparam \Selector28~1 .lut_mask = 64'h777FFFFF777FFFFF;
defparam \Selector28~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_2),
	.datac(!ctrl_opcode_0),
	.datad(!\Selector9~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h0004000400040004;
defparam \Selector25~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~1 (
	.dataa(!logical_ch_addr[3]),
	.datab(!\Selector2~0_combout ),
	.datac(!\Selector7~1_combout ),
	.datad(!ctrl_addr_3),
	.datae(!\Selector25~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~1 .extended_lut = "off";
defparam \Selector25~1 .lut_mask = 64'hEEE00000EEE00000;
defparam \Selector25~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~2 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_3),
	.datac(!\Selector27~0_combout ),
	.datad(!\Selector25~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~2 .extended_lut = "off";
defparam \Selector25~2 .lut_mask = 64'hFF1FFF1FFF1FFF1F;
defparam \Selector25~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~1 (
	.dataa(!ctrl_lock),
	.datab(!\Selector4~0_combout ),
	.datac(!\Selector12~2_combout ),
	.datad(!\WideOr17~0_combout ),
	.datae(!\Selector16~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~1 .extended_lut = "off";
defparam \Selector16~1 .lut_mask = 64'hFFFFFF3BFFFFFF3B;
defparam \Selector16~1 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[5]~0 (
	.dataa(!\Selector3~9_combout ),
	.datab(!\Selector3~7_combout ),
	.datac(!\Selector3~10_combout ),
	.datad(!\WideOr2~combout ),
	.datae(!\Selector3~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[5]~0 .extended_lut = "off";
defparam \master_writedata[5]~0 .lut_mask = 64'h0002000000020000;
defparam \master_writedata[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[5]~1 (
	.dataa(!\Selector3~15_combout ),
	.datab(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datac(!\Selector3~10_combout ),
	.datad(!\Selector3~14_combout ),
	.datae(!\Selector7~1_combout ),
	.dataf(!\master_writedata[5]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[5]~1 .extended_lut = "off";
defparam \master_writedata[5]~1 .lut_mask = 64'hFFFD0000555D0000;
defparam \master_writedata[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[5]~2 (
	.dataa(!\Selector2~0_combout ),
	.datab(!\Selector8~1_combout ),
	.datac(!\Selector7~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[5]~2 .extended_lut = "off";
defparam \master_writedata[5]~2 .lut_mask = 64'h8C8C8C8C8C8C8C8C;
defparam \master_writedata[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!logical_ch_addr[4]),
	.datab(!ctrl_addr_4),
	.datac(!\master_writedata[5]~1_combout ),
	.datad(!\master_writedata[5]~2_combout ),
	.datae(!ctrl_wdata_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h0530F5300530F530;
defparam \Selector24~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector23~0 (
	.dataa(!logical_ch_addr[5]),
	.datab(!\master_writedata[5]~1_combout ),
	.datac(!\master_writedata[5]~2_combout ),
	.datad(!ctrl_addr_5),
	.datae(!ctrl_wdata_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h101CD0DC101CD0DC;
defparam \Selector23~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector22~0 (
	.dataa(!logical_ch_addr[6]),
	.datab(!\master_writedata[5]~1_combout ),
	.datac(!\master_writedata[5]~2_combout ),
	.datad(!ctrl_addr_6),
	.datae(!ctrl_wdata_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector22~0 .extended_lut = "off";
defparam \Selector22~0 .lut_mask = 64'h101CD0DC101CD0DC;
defparam \Selector22~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector21~0 (
	.dataa(!logical_ch_addr[7]),
	.datab(!\master_writedata[5]~1_combout ),
	.datac(!\master_writedata[5]~2_combout ),
	.datad(!ctrl_addr_7),
	.datae(!ctrl_wdata_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~0 .extended_lut = "off";
defparam \Selector21~0 .lut_mask = 64'h101CD0DC101CD0DC;
defparam \Selector21~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!logical_ch_addr[8]),
	.datab(!\master_writedata[5]~1_combout ),
	.datac(!\master_writedata[5]~2_combout ),
	.datad(!ctrl_addr_8),
	.datae(!ctrl_wdata_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h101CD0DC101CD0DC;
defparam \Selector20~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!logical_ch_addr[9]),
	.datab(!\master_writedata[5]~1_combout ),
	.datac(!\master_writedata[5]~2_combout ),
	.datad(!ctrl_addr_9),
	.datae(!ctrl_wdata_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h101CD0DC101CD0DC;
defparam \Selector19~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!\Selector8~1_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(!ctrl_wdata_10),
	.datad(!ctrl_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h0537053705370537;
defparam \Selector18~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!\Selector8~1_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(!ctrl_wdata_11),
	.datad(!ctrl_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'h0537053705370537;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~3 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~3 .extended_lut = "off";
defparam \master_writedata~3 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~3 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~4 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~4 .extended_lut = "off";
defparam \master_writedata~4 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~4 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~5 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~5 .extended_lut = "off";
defparam \master_writedata~5 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~5 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~6 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~6 .extended_lut = "off";
defparam \master_writedata~6 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~6 .shared_arith = "off";

cyclonev_lcell_comb \readdata_for_user[0]~0 (
	.dataa(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.datab(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datac(!\Selector12~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata_for_user[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata_for_user[0]~0 .extended_lut = "off";
defparam \readdata_for_user[0]~0 .lut_mask = 64'h0707070707070707;
defparam \readdata_for_user[0]~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_uif_1 (
	user_reconfig_readdata_12,
	user_reconfig_readdata_13,
	user_reconfig_readdata_14,
	user_reconfig_readdata_15,
	user_reconfig_readdata_16,
	user_reconfig_readdata_17,
	user_reconfig_readdata_18,
	user_reconfig_readdata_19,
	user_reconfig_readdata_20,
	user_reconfig_readdata_21,
	user_reconfig_readdata_22,
	user_reconfig_readdata_23,
	user_reconfig_readdata_24,
	user_reconfig_readdata_25,
	user_reconfig_readdata_26,
	user_reconfig_readdata_27,
	user_reconfig_readdata_28,
	user_reconfig_readdata_29,
	user_reconfig_readdata_30,
	user_reconfig_readdata_31,
	uif_rdata_5,
	uif_rdata_6,
	uif_rdata_7,
	uif_rdata_8,
	uif_rdata_9,
	uif_rdata_10,
	uif_rdata_11,
	uif_rdata_12,
	uif_rdata_13,
	uif_rdata_14,
	uif_rdata_15,
	uif_rdata_16,
	uif_rdata_17,
	uif_rdata_18,
	uif_rdata_19,
	uif_rdata_20,
	uif_rdata_21,
	uif_rdata_22,
	uif_rdata_23,
	uif_rdata_24,
	uif_rdata_25,
	uif_rdata_26,
	uif_rdata_27,
	uif_rdata_28,
	uif_rdata_29,
	uif_rdata_30,
	uif_rdata_31,
	user_reconfig_readdata_0,
	Equal3,
	user_reconfig_readdata_1,
	user_reconfig_readdata_2,
	user_reconfig_readdata_3,
	user_reconfig_readdata_4,
	user_reconfig_readdata_5,
	user_reconfig_readdata_6,
	user_reconfig_readdata_7,
	reconfig_mgmt_readdata_8,
	user_reconfig_readdata_8,
	user_reconfig_readdata_9,
	user_reconfig_readdata_10,
	user_reconfig_readdata_11,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	uif_busy,
	ifsel_notdone_resync,
	uif_writedata_0,
	uif_mode_1,
	uif_mode_0,
	Equal5,
	uif_rdata_0,
	ph_readdata_0,
	uif_logical_ch_addr_0,
	uif_addr_offset_0,
	comb,
	uif_writedata_1,
	uif_rdata_1,
	ph_readdata_1,
	uif_logical_ch_addr_1,
	uif_addr_offset_1,
	uif_writedata_2,
	uif_logical_ch_addr_2,
	ph_readdata_2,
	uif_ctrl_0,
	uif_addr_offset_2,
	uif_rdata_2,
	uif_writedata_3,
	uif_logical_ch_addr_3,
	ph_readdata_3,
	uif_ctrl_1,
	uif_addr_offset_3,
	uif_rdata_3,
	user_reconfig_readdata_101,
	uif_writedata_4,
	uif_rdata_4,
	ph_readdata_4,
	uif_logical_ch_addr_4,
	uif_addr_offset_4,
	uif_writedata_5,
	ph_readdata_5,
	uif_logical_ch_addr_5,
	uif_addr_offset_5,
	uif_writedata_6,
	ph_readdata_6,
	uif_logical_ch_addr_6,
	uif_addr_offset_6,
	uif_writedata_7,
	ph_readdata_7,
	uif_logical_ch_addr_7,
	uif_addr_offset_7,
	uif_writedata_8,
	uif_logical_ch_addr_8,
	ph_readdata_8,
	uif_addr_offset_8,
	uif_writedata_9,
	uif_logical_ch_addr_9,
	ph_readdata_9,
	uif_addr_err,
	illegal_phy_ch,
	uif_addr_offset_9,
	ph_readdata_10,
	uif_writedata_10,
	uif_addr_offset_10,
	ph_readdata_11,
	uif_writedata_11,
	uif_addr_offset_11,
	ph_readdata_12,
	uif_writedata_12,
	ph_readdata_13,
	uif_writedata_13,
	ph_readdata_14,
	uif_writedata_14,
	ph_readdata_15,
	uif_writedata_15,
	ph_readdata_16,
	uif_writedata_16,
	ph_readdata_17,
	uif_writedata_17,
	ph_readdata_18,
	uif_writedata_18,
	ph_readdata_19,
	uif_writedata_19,
	ph_readdata_20,
	uif_writedata_20,
	ph_readdata_21,
	uif_writedata_21,
	ph_readdata_22,
	uif_writedata_22,
	ph_readdata_23,
	uif_writedata_23,
	ph_readdata_24,
	uif_writedata_24,
	ph_readdata_25,
	uif_writedata_25,
	ph_readdata_26,
	uif_writedata_26,
	ph_readdata_27,
	uif_writedata_27,
	ph_readdata_28,
	uif_writedata_28,
	ph_readdata_29,
	uif_writedata_29,
	ph_readdata_30,
	uif_writedata_30,
	ph_readdata_31,
	uif_writedata_31,
	uif_mode_01,
	Mux0,
	Mux3,
	uif_go1,
	WideOr0,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
output 	user_reconfig_readdata_20;
output 	user_reconfig_readdata_21;
output 	user_reconfig_readdata_22;
output 	user_reconfig_readdata_23;
output 	user_reconfig_readdata_24;
output 	user_reconfig_readdata_25;
output 	user_reconfig_readdata_26;
output 	user_reconfig_readdata_27;
output 	user_reconfig_readdata_28;
output 	user_reconfig_readdata_29;
output 	user_reconfig_readdata_30;
output 	user_reconfig_readdata_31;
input 	uif_rdata_5;
input 	uif_rdata_6;
input 	uif_rdata_7;
input 	uif_rdata_8;
input 	uif_rdata_9;
input 	uif_rdata_10;
input 	uif_rdata_11;
input 	uif_rdata_12;
input 	uif_rdata_13;
input 	uif_rdata_14;
input 	uif_rdata_15;
input 	uif_rdata_16;
input 	uif_rdata_17;
input 	uif_rdata_18;
input 	uif_rdata_19;
input 	uif_rdata_20;
input 	uif_rdata_21;
input 	uif_rdata_22;
input 	uif_rdata_23;
input 	uif_rdata_24;
input 	uif_rdata_25;
input 	uif_rdata_26;
input 	uif_rdata_27;
input 	uif_rdata_28;
input 	uif_rdata_29;
input 	uif_rdata_30;
input 	uif_rdata_31;
output 	user_reconfig_readdata_0;
input 	Equal3;
output 	user_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
output 	user_reconfig_readdata_6;
output 	user_reconfig_readdata_7;
input 	reconfig_mgmt_readdata_8;
output 	user_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
output 	user_reconfig_readdata_10;
output 	user_reconfig_readdata_11;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
input 	uif_busy;
input 	ifsel_notdone_resync;
output 	uif_writedata_0;
output 	uif_mode_1;
output 	uif_mode_0;
input 	Equal5;
input 	uif_rdata_0;
input 	ph_readdata_0;
output 	uif_logical_ch_addr_0;
output 	uif_addr_offset_0;
input 	comb;
output 	uif_writedata_1;
input 	uif_rdata_1;
input 	ph_readdata_1;
output 	uif_logical_ch_addr_1;
output 	uif_addr_offset_1;
output 	uif_writedata_2;
output 	uif_logical_ch_addr_2;
input 	ph_readdata_2;
output 	uif_ctrl_0;
output 	uif_addr_offset_2;
input 	uif_rdata_2;
output 	uif_writedata_3;
output 	uif_logical_ch_addr_3;
input 	ph_readdata_3;
output 	uif_ctrl_1;
output 	uif_addr_offset_3;
input 	uif_rdata_3;
input 	user_reconfig_readdata_101;
output 	uif_writedata_4;
input 	uif_rdata_4;
input 	ph_readdata_4;
output 	uif_logical_ch_addr_4;
output 	uif_addr_offset_4;
output 	uif_writedata_5;
input 	ph_readdata_5;
output 	uif_logical_ch_addr_5;
output 	uif_addr_offset_5;
output 	uif_writedata_6;
input 	ph_readdata_6;
output 	uif_logical_ch_addr_6;
output 	uif_addr_offset_6;
output 	uif_writedata_7;
input 	ph_readdata_7;
output 	uif_logical_ch_addr_7;
output 	uif_addr_offset_7;
output 	uif_writedata_8;
output 	uif_logical_ch_addr_8;
input 	ph_readdata_8;
output 	uif_addr_offset_8;
output 	uif_writedata_9;
output 	uif_logical_ch_addr_9;
input 	ph_readdata_9;
input 	uif_addr_err;
input 	illegal_phy_ch;
output 	uif_addr_offset_9;
input 	ph_readdata_10;
output 	uif_writedata_10;
output 	uif_addr_offset_10;
input 	ph_readdata_11;
output 	uif_writedata_11;
output 	uif_addr_offset_11;
input 	ph_readdata_12;
output 	uif_writedata_12;
input 	ph_readdata_13;
output 	uif_writedata_13;
input 	ph_readdata_14;
output 	uif_writedata_14;
input 	ph_readdata_15;
output 	uif_writedata_15;
input 	ph_readdata_16;
output 	uif_writedata_16;
input 	ph_readdata_17;
output 	uif_writedata_17;
input 	ph_readdata_18;
output 	uif_writedata_18;
input 	ph_readdata_19;
output 	uif_writedata_19;
input 	ph_readdata_20;
output 	uif_writedata_20;
input 	ph_readdata_21;
output 	uif_writedata_21;
input 	ph_readdata_22;
output 	uif_writedata_22;
input 	ph_readdata_23;
output 	uif_writedata_23;
input 	ph_readdata_24;
output 	uif_writedata_24;
input 	ph_readdata_25;
output 	uif_writedata_25;
input 	ph_readdata_26;
output 	uif_writedata_26;
input 	ph_readdata_27;
output 	uif_writedata_27;
input 	ph_readdata_28;
output 	uif_writedata_28;
input 	ph_readdata_29;
output 	uif_writedata_29;
input 	ph_readdata_30;
output 	uif_writedata_30;
input 	ph_readdata_31;
output 	uif_writedata_31;
input 	uif_mode_01;
input 	Mux0;
input 	Mux3;
output 	uif_go1;
input 	WideOr0;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux23~0_combout ;
wire \user_reconfig_readdata[10]~6_combout ;
wire \Mux22~0_combout ;
wire \Mux21~0_combout ;
wire \Mux20~0_combout ;
wire \Mux19~0_combout ;
wire \Mux18~0_combout ;
wire \Mux17~0_combout ;
wire \Mux16~0_combout ;
wire \Mux15~0_combout ;
wire \Mux14~0_combout ;
wire \Mux13~0_combout ;
wire \Mux12~0_combout ;
wire \Mux11~0_combout ;
wire \Mux10~0_combout ;
wire \Mux9~0_combout ;
wire \Mux8~0_combout ;
wire \Mux7~0_combout ;
wire \Mux6~0_combout ;
wire \Mux5~0_combout ;
wire \Mux4~0_combout ;
wire \user_reconfig_readdata[0]~0_combout ;
wire \user_reconfig_readdata[0]~1_combout ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \user_reconfig_readdata[0]~2_combout ;
wire \user_reconfig_readdata[0]~3_combout ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \illegal_addr_error~0_combout ;
wire \illegal_addr_error~q ;
wire \int_status_error~combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \user_reconfig_readdata[11]~4_combout ;
wire \user_reconfig_readdata[11]~5_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \always0~0_combout ;
wire \uif_writedata[0]~0_combout ;
wire \uif_mode[1]~1_combout ;
wire \Mux0~0_combout ;
wire \uif_mode[2]~0_combout ;
wire \uif_logical_ch_addr[0]~0_combout ;
wire \uif_addr_offset[0]~0_combout ;
wire \uif_ctrl[1]~0_combout ;
wire \Mux0~1_combout ;


RECONFIGURE_IP_altera_wait_generate_1 wait_gen(
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg1(launch_reg),
	.wait_reg1(wait_reg),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.launch_signal(comb),
	.mgmt_clk_clk(mgmt_clk_clk));

dffeas \user_reconfig_readdata[12] (
	.clk(mgmt_clk_clk),
	.d(\Mux23~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_12),
	.prn(vcc));
defparam \user_reconfig_readdata[12] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[12] .power_up = "low";

dffeas \user_reconfig_readdata[13] (
	.clk(mgmt_clk_clk),
	.d(\Mux22~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_13),
	.prn(vcc));
defparam \user_reconfig_readdata[13] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[13] .power_up = "low";

dffeas \user_reconfig_readdata[14] (
	.clk(mgmt_clk_clk),
	.d(\Mux21~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_14),
	.prn(vcc));
defparam \user_reconfig_readdata[14] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[14] .power_up = "low";

dffeas \user_reconfig_readdata[15] (
	.clk(mgmt_clk_clk),
	.d(\Mux20~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_15),
	.prn(vcc));
defparam \user_reconfig_readdata[15] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[15] .power_up = "low";

dffeas \user_reconfig_readdata[16] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_16),
	.prn(vcc));
defparam \user_reconfig_readdata[16] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[16] .power_up = "low";

dffeas \user_reconfig_readdata[17] (
	.clk(mgmt_clk_clk),
	.d(\Mux18~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_17),
	.prn(vcc));
defparam \user_reconfig_readdata[17] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[17] .power_up = "low";

dffeas \user_reconfig_readdata[18] (
	.clk(mgmt_clk_clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_18),
	.prn(vcc));
defparam \user_reconfig_readdata[18] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[18] .power_up = "low";

dffeas \user_reconfig_readdata[19] (
	.clk(mgmt_clk_clk),
	.d(\Mux16~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_19),
	.prn(vcc));
defparam \user_reconfig_readdata[19] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[19] .power_up = "low";

dffeas \user_reconfig_readdata[20] (
	.clk(mgmt_clk_clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_20),
	.prn(vcc));
defparam \user_reconfig_readdata[20] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[20] .power_up = "low";

dffeas \user_reconfig_readdata[21] (
	.clk(mgmt_clk_clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_21),
	.prn(vcc));
defparam \user_reconfig_readdata[21] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[21] .power_up = "low";

dffeas \user_reconfig_readdata[22] (
	.clk(mgmt_clk_clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_22),
	.prn(vcc));
defparam \user_reconfig_readdata[22] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[22] .power_up = "low";

dffeas \user_reconfig_readdata[23] (
	.clk(mgmt_clk_clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_23),
	.prn(vcc));
defparam \user_reconfig_readdata[23] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[23] .power_up = "low";

dffeas \user_reconfig_readdata[24] (
	.clk(mgmt_clk_clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_24),
	.prn(vcc));
defparam \user_reconfig_readdata[24] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[24] .power_up = "low";

dffeas \user_reconfig_readdata[25] (
	.clk(mgmt_clk_clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_25),
	.prn(vcc));
defparam \user_reconfig_readdata[25] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[25] .power_up = "low";

dffeas \user_reconfig_readdata[26] (
	.clk(mgmt_clk_clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_26),
	.prn(vcc));
defparam \user_reconfig_readdata[26] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[26] .power_up = "low";

dffeas \user_reconfig_readdata[27] (
	.clk(mgmt_clk_clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_27),
	.prn(vcc));
defparam \user_reconfig_readdata[27] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[27] .power_up = "low";

dffeas \user_reconfig_readdata[28] (
	.clk(mgmt_clk_clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_28),
	.prn(vcc));
defparam \user_reconfig_readdata[28] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[28] .power_up = "low";

dffeas \user_reconfig_readdata[29] (
	.clk(mgmt_clk_clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_29),
	.prn(vcc));
defparam \user_reconfig_readdata[29] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[29] .power_up = "low";

dffeas \user_reconfig_readdata[30] (
	.clk(mgmt_clk_clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_30),
	.prn(vcc));
defparam \user_reconfig_readdata[30] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[30] .power_up = "low";

dffeas \user_reconfig_readdata[31] (
	.clk(mgmt_clk_clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_31),
	.prn(vcc));
defparam \user_reconfig_readdata[31] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[31] .power_up = "low";

dffeas \user_reconfig_readdata[0] (
	.clk(mgmt_clk_clk),
	.d(\Mux35~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_0),
	.prn(vcc));
defparam \user_reconfig_readdata[0] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[0] .power_up = "low";

dffeas \user_reconfig_readdata[1] (
	.clk(mgmt_clk_clk),
	.d(\Mux34~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_1),
	.prn(vcc));
defparam \user_reconfig_readdata[1] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[1] .power_up = "low";

dffeas \user_reconfig_readdata[2] (
	.clk(mgmt_clk_clk),
	.d(\Mux33~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_2),
	.prn(vcc));
defparam \user_reconfig_readdata[2] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[2] .power_up = "low";

dffeas \user_reconfig_readdata[3] (
	.clk(mgmt_clk_clk),
	.d(\Mux32~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_3),
	.prn(vcc));
defparam \user_reconfig_readdata[3] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[3] .power_up = "low";

dffeas \user_reconfig_readdata[4] (
	.clk(mgmt_clk_clk),
	.d(\Mux31~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_4),
	.prn(vcc));
defparam \user_reconfig_readdata[4] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[4] .power_up = "low";

dffeas \user_reconfig_readdata[5] (
	.clk(mgmt_clk_clk),
	.d(\Mux30~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_5),
	.prn(vcc));
defparam \user_reconfig_readdata[5] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[5] .power_up = "low";

dffeas \user_reconfig_readdata[6] (
	.clk(mgmt_clk_clk),
	.d(\Mux29~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_6),
	.prn(vcc));
defparam \user_reconfig_readdata[6] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[6] .power_up = "low";

dffeas \user_reconfig_readdata[7] (
	.clk(mgmt_clk_clk),
	.d(\Mux28~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_7),
	.prn(vcc));
defparam \user_reconfig_readdata[7] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[7] .power_up = "low";

dffeas \user_reconfig_readdata[8] (
	.clk(mgmt_clk_clk),
	.d(\Mux27~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_8),
	.prn(vcc));
defparam \user_reconfig_readdata[8] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[8] .power_up = "low";

dffeas \user_reconfig_readdata[9] (
	.clk(mgmt_clk_clk),
	.d(\Mux26~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_9),
	.prn(vcc));
defparam \user_reconfig_readdata[9] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[9] .power_up = "low";

dffeas \user_reconfig_readdata[10] (
	.clk(mgmt_clk_clk),
	.d(\Mux25~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_10),
	.prn(vcc));
defparam \user_reconfig_readdata[10] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[10] .power_up = "low";

dffeas \user_reconfig_readdata[11] (
	.clk(mgmt_clk_clk),
	.d(\Mux24~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[10]~6_combout ),
	.q(user_reconfig_readdata_11),
	.prn(vcc));
defparam \user_reconfig_readdata[11] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[11] .power_up = "low";

dffeas \uif_writedata[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_0),
	.prn(vcc));
defparam \uif_writedata[0] .is_wysiwyg = "true";
defparam \uif_writedata[0] .power_up = "low";

dffeas \uif_mode[1] (
	.clk(mgmt_clk_clk),
	.d(\uif_mode[1]~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_mode[2]~0_combout ),
	.q(uif_mode_1),
	.prn(vcc));
defparam \uif_mode[1] .is_wysiwyg = "true";
defparam \uif_mode[1] .power_up = "low";

dffeas \uif_mode[0] (
	.clk(mgmt_clk_clk),
	.d(Mux3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_mode[2]~0_combout ),
	.q(uif_mode_0),
	.prn(vcc));
defparam \uif_mode[0] .is_wysiwyg = "true";
defparam \uif_mode[0] .power_up = "low";

dffeas \uif_logical_ch_addr[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_0),
	.prn(vcc));
defparam \uif_logical_ch_addr[0] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[0] .power_up = "low";

dffeas \uif_addr_offset[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_0),
	.prn(vcc));
defparam \uif_addr_offset[0] .is_wysiwyg = "true";
defparam \uif_addr_offset[0] .power_up = "low";

dffeas \uif_writedata[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_1),
	.prn(vcc));
defparam \uif_writedata[1] .is_wysiwyg = "true";
defparam \uif_writedata[1] .power_up = "low";

dffeas \uif_logical_ch_addr[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_1),
	.prn(vcc));
defparam \uif_logical_ch_addr[1] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[1] .power_up = "low";

dffeas \uif_addr_offset[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_1),
	.prn(vcc));
defparam \uif_addr_offset[1] .is_wysiwyg = "true";
defparam \uif_addr_offset[1] .power_up = "low";

dffeas \uif_writedata[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_2),
	.prn(vcc));
defparam \uif_writedata[2] .is_wysiwyg = "true";
defparam \uif_writedata[2] .power_up = "low";

dffeas \uif_logical_ch_addr[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_2),
	.prn(vcc));
defparam \uif_logical_ch_addr[2] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[2] .power_up = "low";

dffeas \uif_ctrl[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_ctrl[1]~0_combout ),
	.q(uif_ctrl_0),
	.prn(vcc));
defparam \uif_ctrl[0] .is_wysiwyg = "true";
defparam \uif_ctrl[0] .power_up = "low";

dffeas \uif_addr_offset[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_2),
	.prn(vcc));
defparam \uif_addr_offset[2] .is_wysiwyg = "true";
defparam \uif_addr_offset[2] .power_up = "low";

dffeas \uif_writedata[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_3),
	.prn(vcc));
defparam \uif_writedata[3] .is_wysiwyg = "true";
defparam \uif_writedata[3] .power_up = "low";

dffeas \uif_logical_ch_addr[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_3),
	.prn(vcc));
defparam \uif_logical_ch_addr[3] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[3] .power_up = "low";

dffeas \uif_ctrl[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_ctrl[1]~0_combout ),
	.q(uif_ctrl_1),
	.prn(vcc));
defparam \uif_ctrl[1] .is_wysiwyg = "true";
defparam \uif_ctrl[1] .power_up = "low";

dffeas \uif_addr_offset[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_3),
	.prn(vcc));
defparam \uif_addr_offset[3] .is_wysiwyg = "true";
defparam \uif_addr_offset[3] .power_up = "low";

dffeas \uif_writedata[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_4),
	.prn(vcc));
defparam \uif_writedata[4] .is_wysiwyg = "true";
defparam \uif_writedata[4] .power_up = "low";

dffeas \uif_logical_ch_addr[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_4),
	.prn(vcc));
defparam \uif_logical_ch_addr[4] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[4] .power_up = "low";

dffeas \uif_addr_offset[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_4),
	.prn(vcc));
defparam \uif_addr_offset[4] .is_wysiwyg = "true";
defparam \uif_addr_offset[4] .power_up = "low";

dffeas \uif_writedata[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_5),
	.prn(vcc));
defparam \uif_writedata[5] .is_wysiwyg = "true";
defparam \uif_writedata[5] .power_up = "low";

dffeas \uif_logical_ch_addr[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_5),
	.prn(vcc));
defparam \uif_logical_ch_addr[5] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[5] .power_up = "low";

dffeas \uif_addr_offset[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_5),
	.prn(vcc));
defparam \uif_addr_offset[5] .is_wysiwyg = "true";
defparam \uif_addr_offset[5] .power_up = "low";

dffeas \uif_writedata[6] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_6),
	.prn(vcc));
defparam \uif_writedata[6] .is_wysiwyg = "true";
defparam \uif_writedata[6] .power_up = "low";

dffeas \uif_logical_ch_addr[6] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_6),
	.prn(vcc));
defparam \uif_logical_ch_addr[6] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[6] .power_up = "low";

dffeas \uif_addr_offset[6] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_6),
	.prn(vcc));
defparam \uif_addr_offset[6] .is_wysiwyg = "true";
defparam \uif_addr_offset[6] .power_up = "low";

dffeas \uif_writedata[7] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_7),
	.prn(vcc));
defparam \uif_writedata[7] .is_wysiwyg = "true";
defparam \uif_writedata[7] .power_up = "low";

dffeas \uif_logical_ch_addr[7] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_7),
	.prn(vcc));
defparam \uif_logical_ch_addr[7] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[7] .power_up = "low";

dffeas \uif_addr_offset[7] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_7),
	.prn(vcc));
defparam \uif_addr_offset[7] .is_wysiwyg = "true";
defparam \uif_addr_offset[7] .power_up = "low";

dffeas \uif_writedata[8] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_8),
	.prn(vcc));
defparam \uif_writedata[8] .is_wysiwyg = "true";
defparam \uif_writedata[8] .power_up = "low";

dffeas \uif_logical_ch_addr[8] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_8),
	.prn(vcc));
defparam \uif_logical_ch_addr[8] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[8] .power_up = "low";

dffeas \uif_addr_offset[8] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_8),
	.prn(vcc));
defparam \uif_addr_offset[8] .is_wysiwyg = "true";
defparam \uif_addr_offset[8] .power_up = "low";

dffeas \uif_writedata[9] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_9),
	.prn(vcc));
defparam \uif_writedata[9] .is_wysiwyg = "true";
defparam \uif_writedata[9] .power_up = "low";

dffeas \uif_logical_ch_addr[9] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_9),
	.prn(vcc));
defparam \uif_logical_ch_addr[9] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[9] .power_up = "low";

dffeas \uif_addr_offset[9] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_9),
	.prn(vcc));
defparam \uif_addr_offset[9] .is_wysiwyg = "true";
defparam \uif_addr_offset[9] .power_up = "low";

dffeas \uif_writedata[10] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_10),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_10),
	.prn(vcc));
defparam \uif_writedata[10] .is_wysiwyg = "true";
defparam \uif_writedata[10] .power_up = "low";

dffeas \uif_addr_offset[10] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_10),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_10),
	.prn(vcc));
defparam \uif_addr_offset[10] .is_wysiwyg = "true";
defparam \uif_addr_offset[10] .power_up = "low";

dffeas \uif_writedata[11] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_11),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_11),
	.prn(vcc));
defparam \uif_writedata[11] .is_wysiwyg = "true";
defparam \uif_writedata[11] .power_up = "low";

dffeas \uif_addr_offset[11] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_11),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[0]~0_combout ),
	.q(uif_addr_offset_11),
	.prn(vcc));
defparam \uif_addr_offset[11] .is_wysiwyg = "true";
defparam \uif_addr_offset[11] .power_up = "low";

dffeas \uif_writedata[12] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_12),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_12),
	.prn(vcc));
defparam \uif_writedata[12] .is_wysiwyg = "true";
defparam \uif_writedata[12] .power_up = "low";

dffeas \uif_writedata[13] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_13),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_13),
	.prn(vcc));
defparam \uif_writedata[13] .is_wysiwyg = "true";
defparam \uif_writedata[13] .power_up = "low";

dffeas \uif_writedata[14] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_14),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_14),
	.prn(vcc));
defparam \uif_writedata[14] .is_wysiwyg = "true";
defparam \uif_writedata[14] .power_up = "low";

dffeas \uif_writedata[15] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_15),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_15),
	.prn(vcc));
defparam \uif_writedata[15] .is_wysiwyg = "true";
defparam \uif_writedata[15] .power_up = "low";

dffeas \uif_writedata[16] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_16),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_16),
	.prn(vcc));
defparam \uif_writedata[16] .is_wysiwyg = "true";
defparam \uif_writedata[16] .power_up = "low";

dffeas \uif_writedata[17] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_17),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_17),
	.prn(vcc));
defparam \uif_writedata[17] .is_wysiwyg = "true";
defparam \uif_writedata[17] .power_up = "low";

dffeas \uif_writedata[18] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_18),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_18),
	.prn(vcc));
defparam \uif_writedata[18] .is_wysiwyg = "true";
defparam \uif_writedata[18] .power_up = "low";

dffeas \uif_writedata[19] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_19),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_19),
	.prn(vcc));
defparam \uif_writedata[19] .is_wysiwyg = "true";
defparam \uif_writedata[19] .power_up = "low";

dffeas \uif_writedata[20] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_20),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_20),
	.prn(vcc));
defparam \uif_writedata[20] .is_wysiwyg = "true";
defparam \uif_writedata[20] .power_up = "low";

dffeas \uif_writedata[21] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_21),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_21),
	.prn(vcc));
defparam \uif_writedata[21] .is_wysiwyg = "true";
defparam \uif_writedata[21] .power_up = "low";

dffeas \uif_writedata[22] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_22),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_22),
	.prn(vcc));
defparam \uif_writedata[22] .is_wysiwyg = "true";
defparam \uif_writedata[22] .power_up = "low";

dffeas \uif_writedata[23] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_23),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_23),
	.prn(vcc));
defparam \uif_writedata[23] .is_wysiwyg = "true";
defparam \uif_writedata[23] .power_up = "low";

dffeas \uif_writedata[24] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_24),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_24),
	.prn(vcc));
defparam \uif_writedata[24] .is_wysiwyg = "true";
defparam \uif_writedata[24] .power_up = "low";

dffeas \uif_writedata[25] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_25),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_25),
	.prn(vcc));
defparam \uif_writedata[25] .is_wysiwyg = "true";
defparam \uif_writedata[25] .power_up = "low";

dffeas \uif_writedata[26] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_26),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_26),
	.prn(vcc));
defparam \uif_writedata[26] .is_wysiwyg = "true";
defparam \uif_writedata[26] .power_up = "low";

dffeas \uif_writedata[27] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_27),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_27),
	.prn(vcc));
defparam \uif_writedata[27] .is_wysiwyg = "true";
defparam \uif_writedata[27] .power_up = "low";

dffeas \uif_writedata[28] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_28),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_28),
	.prn(vcc));
defparam \uif_writedata[28] .is_wysiwyg = "true";
defparam \uif_writedata[28] .power_up = "low";

dffeas \uif_writedata[29] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_29),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_29),
	.prn(vcc));
defparam \uif_writedata[29] .is_wysiwyg = "true";
defparam \uif_writedata[29] .power_up = "low";

dffeas \uif_writedata[30] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_30),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_30),
	.prn(vcc));
defparam \uif_writedata[30] .is_wysiwyg = "true";
defparam \uif_writedata[30] .power_up = "low";

dffeas \uif_writedata[31] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_31),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_31),
	.prn(vcc));
defparam \uif_writedata[31] .is_wysiwyg = "true";
defparam \uif_writedata[31] .power_up = "low";

dffeas uif_go(
	.clk(mgmt_clk_clk),
	.d(\Mux0~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_go1),
	.prn(vcc));
defparam uif_go.is_wysiwyg = "true";
defparam uif_go.power_up = "low";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_12),
	.datad(!uif_writedata_12),
	.datae(!uif_rdata_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "off";
defparam \Mux23~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux23~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[10]~6 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!comb),
	.datac(!uif_busy),
	.datad(!uif_mode_1),
	.datae(!uif_mode_0),
	.dataf(!user_reconfig_readdata_101),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[10]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[10]~6 .extended_lut = "off";
defparam \user_reconfig_readdata[10]~6 .lut_mask = 64'h3030302033333333;
defparam \user_reconfig_readdata[10]~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_13),
	.datad(!uif_writedata_13),
	.datae(!uif_rdata_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "off";
defparam \Mux22~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux22~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_14),
	.datad(!uif_writedata_14),
	.datae(!uif_rdata_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "off";
defparam \Mux21~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux21~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_15),
	.datad(!uif_writedata_15),
	.datae(!uif_rdata_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "off";
defparam \Mux20~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux20~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_16),
	.datad(!uif_writedata_16),
	.datae(!uif_rdata_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "off";
defparam \Mux19~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_17),
	.datad(!uif_writedata_17),
	.datae(!uif_rdata_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "off";
defparam \Mux18~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux18~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_18),
	.datad(!uif_writedata_18),
	.datae(!uif_rdata_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "off";
defparam \Mux17~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux17~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_19),
	.datad(!uif_writedata_19),
	.datae(!uif_rdata_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "off";
defparam \Mux16~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux16~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_20),
	.datad(!uif_writedata_20),
	.datae(!uif_rdata_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~0 .extended_lut = "off";
defparam \Mux15~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux15~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_21),
	.datad(!uif_writedata_21),
	.datae(!uif_rdata_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "off";
defparam \Mux14~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux14~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_22),
	.datad(!uif_writedata_22),
	.datae(!uif_rdata_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "off";
defparam \Mux13~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux13~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_23),
	.datad(!uif_writedata_23),
	.datae(!uif_rdata_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "off";
defparam \Mux12~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux12~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_24),
	.datad(!uif_writedata_24),
	.datae(!uif_rdata_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "off";
defparam \Mux11~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_25),
	.datad(!uif_writedata_25),
	.datae(!uif_rdata_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_26),
	.datad(!uif_writedata_26),
	.datae(!uif_rdata_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_27),
	.datad(!uif_writedata_27),
	.datae(!uif_rdata_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_28),
	.datad(!uif_writedata_28),
	.datae(!uif_rdata_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_29),
	.datad(!uif_writedata_29),
	.datae(!uif_rdata_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux6~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_30),
	.datad(!uif_writedata_30),
	.datae(!uif_rdata_30),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux5~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal5),
	.datac(!ph_readdata_31),
	.datad(!uif_writedata_31),
	.datae(!uif_rdata_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~0 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~0 .lut_mask = 64'h070F070F070F070F;
defparam \user_reconfig_readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~1 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~1 .lut_mask = 64'h0F070F070F070F07;
defparam \user_reconfig_readdata[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_0),
	.datad(!uif_logical_ch_addr_0),
	.datae(!uif_addr_offset_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~0 .extended_lut = "off";
defparam \Mux35~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux35~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~1 (
	.dataa(!uif_writedata_0),
	.datab(!\user_reconfig_readdata[0]~0_combout ),
	.datac(!\user_reconfig_readdata[0]~1_combout ),
	.datad(!uif_rdata_0),
	.datae(!\Mux35~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux35~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~1 .extended_lut = "off";
defparam \Mux35~1 .lut_mask = 64'h101CD0DC101CD0DC;
defparam \Mux35~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~2 (
	.dataa(!reconfig_mgmt_address_0),
	.datab(!uif_busy),
	.datac(!uif_mode_1),
	.datad(!uif_mode_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~2 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~2 .lut_mask = 64'hCCC4CCC4CCC4CCC4;
defparam \user_reconfig_readdata[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~3 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!comb),
	.datae(!\user_reconfig_readdata[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~3 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~3 .lut_mask = 64'h00D700FF00D700FF;
defparam \user_reconfig_readdata[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_1),
	.datad(!uif_logical_ch_addr_1),
	.datae(!uif_addr_offset_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~0 .extended_lut = "off";
defparam \Mux34~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux34~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_1),
	.datad(!uif_rdata_1),
	.datae(!\Mux34~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux34~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~1 .extended_lut = "off";
defparam \Mux34~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux34~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~0 (
	.dataa(!uif_logical_ch_addr_2),
	.datab(!ph_readdata_2),
	.datac(!uif_ctrl_0),
	.datad(!uif_addr_offset_2),
	.datae(!reconfig_mgmt_address_0),
	.dataf(!reconfig_mgmt_address_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~0 .extended_lut = "off";
defparam \Mux33~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux33~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_2),
	.datad(!\Mux33~0_combout ),
	.datae(!uif_rdata_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux33~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~1 .extended_lut = "off";
defparam \Mux33~1 .lut_mask = 64'h048C26AE048C26AE;
defparam \Mux33~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~0 (
	.dataa(!uif_logical_ch_addr_3),
	.datab(!ph_readdata_3),
	.datac(!uif_ctrl_1),
	.datad(!uif_addr_offset_3),
	.datae(!reconfig_mgmt_address_0),
	.dataf(!reconfig_mgmt_address_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~0 .extended_lut = "off";
defparam \Mux32~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux32~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_3),
	.datad(!\Mux32~0_combout ),
	.datae(!uif_rdata_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~1 .extended_lut = "off";
defparam \Mux32~1 .lut_mask = 64'h048C26AE048C26AE;
defparam \Mux32~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux31~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_4),
	.datad(!uif_logical_ch_addr_4),
	.datae(!uif_addr_offset_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~0 .extended_lut = "off";
defparam \Mux31~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux31~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux31~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_4),
	.datad(!uif_rdata_4),
	.datae(!\Mux31~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux31~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~1 .extended_lut = "off";
defparam \Mux31~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux31~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux30~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_5),
	.datad(!uif_logical_ch_addr_5),
	.datae(!uif_addr_offset_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~0 .extended_lut = "off";
defparam \Mux30~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux30~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux30~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_5),
	.datad(!uif_rdata_5),
	.datae(!\Mux30~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux30~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~1 .extended_lut = "off";
defparam \Mux30~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux30~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux29~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_6),
	.datad(!uif_logical_ch_addr_6),
	.datae(!uif_addr_offset_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~0 .extended_lut = "off";
defparam \Mux29~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux29~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux29~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_6),
	.datad(!uif_rdata_6),
	.datae(!\Mux29~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux29~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~1 .extended_lut = "off";
defparam \Mux29~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux29~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_7),
	.datad(!uif_logical_ch_addr_7),
	.datae(!uif_addr_offset_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~0 .extended_lut = "off";
defparam \Mux28~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux28~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_7),
	.datad(!uif_rdata_7),
	.datae(!\Mux28~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~1 .extended_lut = "off";
defparam \Mux28~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux28~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!uif_logical_ch_addr_8),
	.datab(!ph_readdata_8),
	.datac(!uif_busy),
	.datad(!uif_addr_offset_8),
	.datae(!reconfig_mgmt_address_0),
	.dataf(!reconfig_mgmt_address_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "off";
defparam \Mux27~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_8),
	.datad(!\Mux27~0_combout ),
	.datae(!uif_rdata_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~1 .extended_lut = "off";
defparam \Mux27~1 .lut_mask = 64'h048C26AE048C26AE;
defparam \Mux27~1 .shared_arith = "off";

cyclonev_lcell_comb \illegal_addr_error~0 (
	.dataa(!Equal3),
	.datab(!reconfig_mgmt_read),
	.datac(!reconfig_mgmt_write),
	.datad(!\illegal_addr_error~q ),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\illegal_addr_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \illegal_addr_error~0 .extended_lut = "off";
defparam \illegal_addr_error~0 .lut_mask = 64'h000015FF000015FF;
defparam \illegal_addr_error~0 .shared_arith = "off";

dffeas illegal_addr_error(
	.clk(mgmt_clk_clk),
	.d(\illegal_addr_error~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\illegal_addr_error~q ),
	.prn(vcc));
defparam illegal_addr_error.is_wysiwyg = "true";
defparam illegal_addr_error.power_up = "low";

cyclonev_lcell_comb int_status_error(
	.dataa(!\illegal_addr_error~q ),
	.datab(!uif_addr_err),
	.datac(!illegal_phy_ch),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_status_error~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam int_status_error.extended_lut = "off";
defparam int_status_error.lut_mask = 64'h8080808080808080;
defparam int_status_error.shared_arith = "off";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!uif_logical_ch_addr_9),
	.datab(!ph_readdata_9),
	.datac(!\int_status_error~combout ),
	.datad(!uif_addr_offset_9),
	.datae(!reconfig_mgmt_address_0),
	.dataf(!reconfig_mgmt_address_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "off";
defparam \Mux26~0 .lut_mask = 64'h55553333F0F000FF;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~1 (
	.dataa(!\user_reconfig_readdata[0]~0_combout ),
	.datab(!\user_reconfig_readdata[0]~1_combout ),
	.datac(!uif_writedata_9),
	.datad(!\Mux26~0_combout ),
	.datae(!uif_rdata_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~1 .extended_lut = "off";
defparam \Mux26~1 .lut_mask = 64'h048C26AE048C26AE;
defparam \Mux26~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[11]~4 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[11]~4 .extended_lut = "off";
defparam \user_reconfig_readdata[11]~4 .lut_mask = 64'h2020202020202020;
defparam \user_reconfig_readdata[11]~4 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[11]~5 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[11]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[11]~5 .extended_lut = "off";
defparam \user_reconfig_readdata[11]~5 .lut_mask = 64'h0008000800080008;
defparam \user_reconfig_readdata[11]~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal5),
	.datae(!uif_rdata_10),
	.dataf(!uif_addr_offset_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "off";
defparam \Mux25~0 .lut_mask = 64'h0000080030303830;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~1 (
	.dataa(!ph_readdata_10),
	.datab(!\user_reconfig_readdata[11]~4_combout ),
	.datac(!uif_writedata_10),
	.datad(!\user_reconfig_readdata[11]~5_combout ),
	.datae(!\Mux25~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~1 .extended_lut = "off";
defparam \Mux25~1 .lut_mask = 64'h111DDDDD111DDDDD;
defparam \Mux25~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal5),
	.datae(!uif_rdata_11),
	.dataf(!uif_addr_offset_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "off";
defparam \Mux24~0 .lut_mask = 64'h0000080030303830;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~1 (
	.dataa(!\user_reconfig_readdata[11]~4_combout ),
	.datab(!\user_reconfig_readdata[11]~5_combout ),
	.datac(!ph_readdata_11),
	.datad(!uif_writedata_11),
	.datae(!\Mux24~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~1 .extended_lut = "off";
defparam \Mux24~1 .lut_mask = 64'h0527AFAF0527AFAF;
defparam \Mux24~1 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!Equal3),
	.datab(!reconfig_mgmt_write),
	.datac(!uif_busy),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h1010101010101010;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_writedata[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_writedata[0]~0 .extended_lut = "off";
defparam \uif_writedata[0]~0 .lut_mask = 64'h0008000800080008;
defparam \uif_writedata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_mode[1]~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_mode[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_mode[1]~1 .extended_lut = "off";
defparam \uif_mode[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \uif_mode[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!comb),
	.datab(!uif_busy),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h4444444444444444;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_mode[2]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!uif_mode_01),
	.datac(!Mux0),
	.datad(!\always0~0_combout ),
	.datae(!\Mux0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_mode[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_mode[2]~0 .extended_lut = "off";
defparam \uif_mode[2]~0 .lut_mask = 64'h00040A0E00040A0E;
defparam \uif_mode[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_logical_ch_addr[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_logical_ch_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_logical_ch_addr[0]~0 .extended_lut = "off";
defparam \uif_logical_ch_addr[0]~0 .lut_mask = 64'h0080008000800080;
defparam \uif_logical_ch_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_addr_offset[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_addr_offset[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_addr_offset[0]~0 .extended_lut = "off";
defparam \uif_addr_offset[0]~0 .lut_mask = 64'h0010001000100010;
defparam \uif_addr_offset[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_ctrl[1]~0 (
	.dataa(!reconfig_mgmt_readdata_8),
	.datab(!\always0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_ctrl[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_ctrl[1]~0 .extended_lut = "off";
defparam \uif_ctrl[1]~0 .lut_mask = 64'h1111111111111111;
defparam \uif_ctrl[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!uif_mode_01),
	.datac(!Mux0),
	.datad(!\always0~0_combout ),
	.datae(!\Mux0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~1 .extended_lut = "off";
defparam \Mux0~1 .lut_mask = 64'h00040A0E00040A0E;
defparam \Mux0~1 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_altera_wait_generate_1 (
	resync_chains0sync_r_1,
	launch_reg1,
	wait_reg1,
	ifsel_notdone_resync,
	launch_signal,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
output 	launch_reg1;
output 	wait_reg1;
input 	ifsel_notdone_resync;
input 	launch_signal;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_reg~0_combout ;


RECONFIGURE_IP_alt_xcvr_resync_1 rst_sync(
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.clk(mgmt_clk_clk));

dffeas launch_reg(
	.clk(mgmt_clk_clk),
	.d(launch_signal),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(launch_reg1),
	.prn(vcc));
defparam launch_reg.is_wysiwyg = "true";
defparam launch_reg.power_up = "low";

dffeas wait_reg(
	.clk(mgmt_clk_clk),
	.d(\wait_reg~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_reg1),
	.prn(vcc));
defparam wait_reg.is_wysiwyg = "true";
defparam wait_reg.power_up = "low";

cyclonev_lcell_comb \wait_reg~0 (
	.dataa(!resync_chains0sync_r_1),
	.datab(!launch_signal),
	.datac(!launch_reg1),
	.datad(!wait_reg1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_reg~0 .extended_lut = "off";
defparam \wait_reg~0 .lut_mask = 64'h0100010001000100;
defparam \wait_reg~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_resync_1 (
	resync_chains0sync_r_1,
	ifsel_notdone_resync,
	clk)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
input 	ifsel_notdone_resync;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \resync_chains[0].sync_r[0]~q ;


dffeas \resync_chains[0].sync_r[1] (
	.clk(clk),
	.d(\resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resync_chains0sync_r_1),
	.prn(vcc));
defparam \resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[1] .power_up = "low";

dffeas \resync_chains[0].sync_r[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[0] .power_up = "low";

endmodule

module RECONFIGURE_IP_av_xcvr_reconfig_mif_avmm (
	stream_address_0,
	stream_address_1,
	stream_address_2,
	stream_address_3,
	stream_address_4,
	stream_address_5,
	stream_address_6,
	stream_address_7,
	stream_address_8,
	stream_address_9,
	stream_address_10,
	stream_address_11,
	stream_address_12,
	stream_address_13,
	stream_address_14,
	stream_address_15,
	stream_address_16,
	stream_address_17,
	stream_address_18,
	stream_address_19,
	stream_address_20,
	stream_address_21,
	stream_address_22,
	stream_address_23,
	stream_address_24,
	stream_address_25,
	stream_address_26,
	stream_address_27,
	stream_address_28,
	stream_address_29,
	stream_address_30,
	stream_address_31,
	av_mif_addr_4,
	av_mif_addr_5,
	av_mif_addr_2,
	av_mif_addr_1,
	av_mif_addr_0,
	av_mif_addr_3,
	av_mif_addr_8,
	av_mif_addr_9,
	av_mif_addr_10,
	av_mif_addr_7,
	av_mif_addr_6,
	stream_read1,
	pll_mif_busy,
	reset,
	av_ctrl_req1,
	ctrl_op_done,
	mif_err_reg_4,
	mif_err_reg_1,
	mif_err_reg_0,
	ctrl_av_go,
	pll_go1,
	mif_base_addr_0,
	mif_base_addr_1,
	mif_base_addr_2,
	mif_base_addr_3,
	mif_base_addr_4,
	mif_base_addr_5,
	mif_base_addr_6,
	mif_base_addr_7,
	mif_base_addr_8,
	mif_base_addr_9,
	mif_base_addr_10,
	mif_base_addr_11,
	mif_base_addr_12,
	mif_base_addr_13,
	mif_base_addr_14,
	mif_base_addr_15,
	mif_base_addr_16,
	mif_base_addr_17,
	mif_base_addr_18,
	mif_base_addr_19,
	mif_base_addr_20,
	mif_base_addr_21,
	mif_base_addr_22,
	mif_base_addr_23,
	mif_base_addr_24,
	mif_base_addr_25,
	mif_base_addr_26,
	mif_base_addr_27,
	mif_base_addr_28,
	mif_base_addr_29,
	mif_base_addr_30,
	mif_base_addr_31,
	av_addr_burst1,
	av_opcode_err1,
	av_done1,
	pll_type1,
	mif_rec_data_1,
	mif_rec_addr_7,
	mif_rec_addr_5,
	mif_rec_addr_6,
	mif_rec_data_2,
	mif_rec_data_0,
	mif_rec_data_3,
	av_mif_type_valid1,
	av_mif_type_1,
	av_mif_type_0,
	mif_rec_data_4,
	mif_rec_data_5,
	mif_rec_data_6,
	mif_rec_data_7,
	mif_rec_data_8,
	mif_rec_data_9,
	mif_rec_data_10,
	mif_rec_data_11,
	mif_rec_data_12,
	mif_rec_data_13,
	mif_rec_data_14,
	mif_rec_data_15,
	mif_addr_mode,
	clk,
	reconfig_mif_waitrequest,
	stream_readdata)/* synthesis synthesis_greybox=0 */;
output 	stream_address_0;
output 	stream_address_1;
output 	stream_address_2;
output 	stream_address_3;
output 	stream_address_4;
output 	stream_address_5;
output 	stream_address_6;
output 	stream_address_7;
output 	stream_address_8;
output 	stream_address_9;
output 	stream_address_10;
output 	stream_address_11;
output 	stream_address_12;
output 	stream_address_13;
output 	stream_address_14;
output 	stream_address_15;
output 	stream_address_16;
output 	stream_address_17;
output 	stream_address_18;
output 	stream_address_19;
output 	stream_address_20;
output 	stream_address_21;
output 	stream_address_22;
output 	stream_address_23;
output 	stream_address_24;
output 	stream_address_25;
output 	stream_address_26;
output 	stream_address_27;
output 	stream_address_28;
output 	stream_address_29;
output 	stream_address_30;
output 	stream_address_31;
output 	av_mif_addr_4;
output 	av_mif_addr_5;
output 	av_mif_addr_2;
output 	av_mif_addr_1;
output 	av_mif_addr_0;
output 	av_mif_addr_3;
output 	av_mif_addr_8;
output 	av_mif_addr_9;
output 	av_mif_addr_10;
output 	av_mif_addr_7;
output 	av_mif_addr_6;
output 	stream_read1;
input 	pll_mif_busy;
input 	reset;
output 	av_ctrl_req1;
input 	ctrl_op_done;
input 	mif_err_reg_4;
input 	mif_err_reg_1;
input 	mif_err_reg_0;
input 	ctrl_av_go;
output 	pll_go1;
input 	mif_base_addr_0;
input 	mif_base_addr_1;
input 	mif_base_addr_2;
input 	mif_base_addr_3;
input 	mif_base_addr_4;
input 	mif_base_addr_5;
input 	mif_base_addr_6;
input 	mif_base_addr_7;
input 	mif_base_addr_8;
input 	mif_base_addr_9;
input 	mif_base_addr_10;
input 	mif_base_addr_11;
input 	mif_base_addr_12;
input 	mif_base_addr_13;
input 	mif_base_addr_14;
input 	mif_base_addr_15;
input 	mif_base_addr_16;
input 	mif_base_addr_17;
input 	mif_base_addr_18;
input 	mif_base_addr_19;
input 	mif_base_addr_20;
input 	mif_base_addr_21;
input 	mif_base_addr_22;
input 	mif_base_addr_23;
input 	mif_base_addr_24;
input 	mif_base_addr_25;
input 	mif_base_addr_26;
input 	mif_base_addr_27;
input 	mif_base_addr_28;
input 	mif_base_addr_29;
input 	mif_base_addr_30;
input 	mif_base_addr_31;
output 	av_addr_burst1;
output 	av_opcode_err1;
output 	av_done1;
output 	pll_type1;
output 	mif_rec_data_1;
output 	mif_rec_addr_7;
output 	mif_rec_addr_5;
output 	mif_rec_addr_6;
output 	mif_rec_data_2;
output 	mif_rec_data_0;
output 	mif_rec_data_3;
output 	av_mif_type_valid1;
output 	av_mif_type_1;
output 	av_mif_type_0;
output 	mif_rec_data_4;
output 	mif_rec_data_5;
output 	mif_rec_data_6;
output 	mif_rec_data_7;
output 	mif_rec_data_8;
output 	mif_rec_data_9;
output 	mif_rec_data_10;
output 	mif_rec_data_11;
output 	mif_rec_data_12;
output 	mif_rec_data_13;
output 	mif_rec_data_14;
output 	mif_rec_data_15;
input 	mif_addr_mode;
input 	clk;
input 	reconfig_mif_waitrequest;
input 	[15:0] stream_readdata;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~1_sumout ;
wire \av_state.AV_DEC_HDR~q ;
wire \mif_rec_len[0]~q ;
wire \mif_rec_len[4]~q ;
wire \mif_rec_len[3]~q ;
wire \mif_rec_len[2]~q ;
wire \mif_rec_len[1]~q ;
wire \Equal2~0_combout ;
wire \mif_len_cnt[1]~7_combout ;
wire \mif_len_cnt[1]~q ;
wire \Selector2~1_combout ;
wire \mif_len_cnt[2]~5_combout ;
wire \mif_len_cnt[2]~6_combout ;
wire \mif_len_cnt[2]~q ;
wire \mif_len_cnt[3]~3_combout ;
wire \mif_len_cnt[3]~4_combout ;
wire \mif_len_cnt[3]~q ;
wire \Add2~0_combout ;
wire \mif_len_cnt[4]~2_combout ;
wire \mif_len_cnt[4]~q ;
wire \Equal0~0_combout ;
wire \mif_rec_addr[1]~q ;
wire \mif_rec_addr[0]~q ;
wire \mif_rec_addr[4]~q ;
wire \mif_rec_addr[3]~q ;
wire \mif_rec_addr[2]~q ;
wire \rec_is_eom~0_combout ;
wire \rec_is_eom~1_combout ;
wire \invalid_rec~0_combout ;
wire \mif_strm_active~0_combout ;
wire \mif_strm_active~q ;
wire \invalid_rec~1_combout ;
wire \Selector4~1_combout ;
wire \Selector4~2_combout ;
wire \av_state.AV_REC_ERR~q ;
wire \Selector0~0_combout ;
wire \av_state.AV_IDLE~q ;
wire \Selector3~3_combout ;
wire \Selector3~4_combout ;
wire \av_state.AV_WF_DONE~q ;
wire \Selector1~2_combout ;
wire \pll_active~0_combout ;
wire \pll_active~q ;
wire \pll_active_dly~q ;
wire \Selector4~0_combout ;
wire \Selector3~2_combout ;
wire \Selector2~2_combout ;
wire \Selector2~3_combout ;
wire \av_state.AV_RD_DATA~q ;
wire \mif_rec_data~0_combout ;
wire \mif_len_cnt[4]~0_combout ;
wire \mif_len_cnt[0]~1_combout ;
wire \mif_len_cnt[0]~q ;
wire \Equal6~0_combout ;
wire \rec_is_som~0_combout ;
wire \Selector1~3_combout ;
wire \Selector1~4_combout ;
wire \Selector1~5_combout ;
wire \Selector1~7_combout ;
wire \av_state.AV_RD_HDR~q ;
wire \av_next_state.AV_DEC_HDR~0_combout ;
wire \mif_next_offset~0_combout ;
wire \mif_next_offset[28]~1_combout ;
wire \mif_next_offset[0]~q ;
wire \Add0~1_sumout ;
wire \Selector1~6_combout ;
wire \stream_address~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \mif_next_offset[1]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \mif_next_offset[2]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \mif_next_offset[3]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \mif_next_offset[4]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \mif_next_offset[5]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add1~22 ;
wire \Add1~25_sumout ;
wire \mif_next_offset[6]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add1~26 ;
wire \Add1~29_sumout ;
wire \mif_next_offset[7]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add1~30 ;
wire \Add1~33_sumout ;
wire \mif_next_offset[8]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add1~34 ;
wire \Add1~37_sumout ;
wire \mif_next_offset[9]~q ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add1~38 ;
wire \Add1~41_sumout ;
wire \mif_next_offset[10]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add1~42 ;
wire \Add1~45_sumout ;
wire \mif_next_offset[11]~q ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add1~46 ;
wire \Add1~49_sumout ;
wire \mif_next_offset[12]~q ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add1~50 ;
wire \Add1~53_sumout ;
wire \mif_next_offset[13]~q ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add1~54 ;
wire \Add1~57_sumout ;
wire \mif_next_offset[14]~q ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add1~58 ;
wire \Add1~61_sumout ;
wire \mif_next_offset[15]~q ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add1~62 ;
wire \Add1~65_sumout ;
wire \mif_next_offset[16]~q ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add1~66 ;
wire \Add1~69_sumout ;
wire \mif_next_offset[17]~q ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add1~70 ;
wire \Add1~73_sumout ;
wire \mif_next_offset[18]~q ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add1~74 ;
wire \Add1~77_sumout ;
wire \mif_next_offset[19]~q ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add1~78 ;
wire \Add1~81_sumout ;
wire \mif_next_offset[20]~q ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add1~82 ;
wire \Add1~85_sumout ;
wire \mif_next_offset[21]~q ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add1~86 ;
wire \Add1~89_sumout ;
wire \mif_next_offset[22]~q ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add1~90 ;
wire \Add1~93_sumout ;
wire \mif_next_offset[23]~q ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add1~94 ;
wire \Add1~97_sumout ;
wire \mif_next_offset[24]~q ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add1~98 ;
wire \Add1~101_sumout ;
wire \mif_next_offset[25]~q ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add1~102 ;
wire \Add1~105_sumout ;
wire \mif_next_offset[26]~q ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add1~106 ;
wire \Add1~109_sumout ;
wire \mif_next_offset[27]~q ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add1~110 ;
wire \Add1~113_sumout ;
wire \mif_next_offset[28]~q ;
wire \Add0~110 ;
wire \Add0~113_sumout ;
wire \Add1~114 ;
wire \Add1~117_sumout ;
wire \mif_next_offset[29]~q ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add1~118 ;
wire \Add1~121_sumout ;
wire \mif_next_offset[30]~q ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add1~122 ;
wire \Add1~125_sumout ;
wire \mif_next_offset[31]~q ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add3~18 ;
wire \Add3~14 ;
wire \Add3~10 ;
wire \Add3~22 ;
wire \Add3~1_sumout ;
wire \av_mif_addr[2]~0_combout ;
wire \av_mif_addr[2]~1_combout ;
wire \av_mif_addr[2]~2_combout ;
wire \av_mif_addr[2]~3_combout ;
wire \Add3~2 ;
wire \Add3~5_sumout ;
wire \Add3~9_sumout ;
wire \Add3~13_sumout ;
wire \Add3~17_sumout ;
wire \Add3~21_sumout ;
wire \Add3~6 ;
wire \Add3~42 ;
wire \Add3~38 ;
wire \Add3~25_sumout ;
wire \mif_rec_addr[8]~q ;
wire \Add3~26 ;
wire \Add3~29_sumout ;
wire \mif_rec_addr[9]~q ;
wire \Add3~30 ;
wire \Add3~33_sumout ;
wire \mif_rec_addr[10]~q ;
wire \Add3~37_sumout ;
wire \Add3~41_sumout ;
wire \stream_read~0_combout ;
wire \av_ctrl_req~0_combout ;
wire \pll_go~0_combout ;
wire \always6~0_combout ;
wire \always6~1_combout ;
wire \always6~2_combout ;
wire \always6~3_combout ;
wire \always6~4_combout ;
wire \always6~5_combout ;
wire \always6~6_combout ;
wire \always6~7_combout ;
wire \always6~8_combout ;
wire \always6~9_combout ;
wire \always6~10_combout ;
wire \always6~11_combout ;
wire \always6~12_combout ;
wire \always6~13_combout ;
wire \first_mif_entry~q ;
wire \av_opcode_err~0_combout ;
wire \av_done~0_combout ;
wire \Equal5~0_combout ;
wire \rec_is_cgb~combout ;
wire \rec_is_type~0_combout ;
wire \av_mif_type~0_combout ;
wire \av_mif_type~1_combout ;


dffeas \stream_address[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_0),
	.prn(vcc));
defparam \stream_address[0] .is_wysiwyg = "true";
defparam \stream_address[0] .power_up = "low";

dffeas \stream_address[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_1),
	.prn(vcc));
defparam \stream_address[1] .is_wysiwyg = "true";
defparam \stream_address[1] .power_up = "low";

dffeas \stream_address[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_2),
	.prn(vcc));
defparam \stream_address[2] .is_wysiwyg = "true";
defparam \stream_address[2] .power_up = "low";

dffeas \stream_address[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_3),
	.prn(vcc));
defparam \stream_address[3] .is_wysiwyg = "true";
defparam \stream_address[3] .power_up = "low";

dffeas \stream_address[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_4),
	.prn(vcc));
defparam \stream_address[4] .is_wysiwyg = "true";
defparam \stream_address[4] .power_up = "low";

dffeas \stream_address[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_5),
	.prn(vcc));
defparam \stream_address[5] .is_wysiwyg = "true";
defparam \stream_address[5] .power_up = "low";

dffeas \stream_address[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_6),
	.prn(vcc));
defparam \stream_address[6] .is_wysiwyg = "true";
defparam \stream_address[6] .power_up = "low";

dffeas \stream_address[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_7),
	.prn(vcc));
defparam \stream_address[7] .is_wysiwyg = "true";
defparam \stream_address[7] .power_up = "low";

dffeas \stream_address[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_8),
	.prn(vcc));
defparam \stream_address[8] .is_wysiwyg = "true";
defparam \stream_address[8] .power_up = "low";

dffeas \stream_address[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_9),
	.prn(vcc));
defparam \stream_address[9] .is_wysiwyg = "true";
defparam \stream_address[9] .power_up = "low";

dffeas \stream_address[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_10),
	.prn(vcc));
defparam \stream_address[10] .is_wysiwyg = "true";
defparam \stream_address[10] .power_up = "low";

dffeas \stream_address[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_11),
	.prn(vcc));
defparam \stream_address[11] .is_wysiwyg = "true";
defparam \stream_address[11] .power_up = "low";

dffeas \stream_address[12] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_12),
	.prn(vcc));
defparam \stream_address[12] .is_wysiwyg = "true";
defparam \stream_address[12] .power_up = "low";

dffeas \stream_address[13] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_13),
	.prn(vcc));
defparam \stream_address[13] .is_wysiwyg = "true";
defparam \stream_address[13] .power_up = "low";

dffeas \stream_address[14] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_14),
	.prn(vcc));
defparam \stream_address[14] .is_wysiwyg = "true";
defparam \stream_address[14] .power_up = "low";

dffeas \stream_address[15] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_15),
	.prn(vcc));
defparam \stream_address[15] .is_wysiwyg = "true";
defparam \stream_address[15] .power_up = "low";

dffeas \stream_address[16] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_16),
	.prn(vcc));
defparam \stream_address[16] .is_wysiwyg = "true";
defparam \stream_address[16] .power_up = "low";

dffeas \stream_address[17] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_17),
	.prn(vcc));
defparam \stream_address[17] .is_wysiwyg = "true";
defparam \stream_address[17] .power_up = "low";

dffeas \stream_address[18] (
	.clk(clk),
	.d(\Add0~73_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_18),
	.prn(vcc));
defparam \stream_address[18] .is_wysiwyg = "true";
defparam \stream_address[18] .power_up = "low";

dffeas \stream_address[19] (
	.clk(clk),
	.d(\Add0~77_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_19),
	.prn(vcc));
defparam \stream_address[19] .is_wysiwyg = "true";
defparam \stream_address[19] .power_up = "low";

dffeas \stream_address[20] (
	.clk(clk),
	.d(\Add0~81_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_20),
	.prn(vcc));
defparam \stream_address[20] .is_wysiwyg = "true";
defparam \stream_address[20] .power_up = "low";

dffeas \stream_address[21] (
	.clk(clk),
	.d(\Add0~85_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_21),
	.prn(vcc));
defparam \stream_address[21] .is_wysiwyg = "true";
defparam \stream_address[21] .power_up = "low";

dffeas \stream_address[22] (
	.clk(clk),
	.d(\Add0~89_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_22),
	.prn(vcc));
defparam \stream_address[22] .is_wysiwyg = "true";
defparam \stream_address[22] .power_up = "low";

dffeas \stream_address[23] (
	.clk(clk),
	.d(\Add0~93_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_23),
	.prn(vcc));
defparam \stream_address[23] .is_wysiwyg = "true";
defparam \stream_address[23] .power_up = "low";

dffeas \stream_address[24] (
	.clk(clk),
	.d(\Add0~97_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_24),
	.prn(vcc));
defparam \stream_address[24] .is_wysiwyg = "true";
defparam \stream_address[24] .power_up = "low";

dffeas \stream_address[25] (
	.clk(clk),
	.d(\Add0~101_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_25),
	.prn(vcc));
defparam \stream_address[25] .is_wysiwyg = "true";
defparam \stream_address[25] .power_up = "low";

dffeas \stream_address[26] (
	.clk(clk),
	.d(\Add0~105_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_26),
	.prn(vcc));
defparam \stream_address[26] .is_wysiwyg = "true";
defparam \stream_address[26] .power_up = "low";

dffeas \stream_address[27] (
	.clk(clk),
	.d(\Add0~109_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_27),
	.prn(vcc));
defparam \stream_address[27] .is_wysiwyg = "true";
defparam \stream_address[27] .power_up = "low";

dffeas \stream_address[28] (
	.clk(clk),
	.d(\Add0~113_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_28),
	.prn(vcc));
defparam \stream_address[28] .is_wysiwyg = "true";
defparam \stream_address[28] .power_up = "low";

dffeas \stream_address[29] (
	.clk(clk),
	.d(\Add0~117_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_29),
	.prn(vcc));
defparam \stream_address[29] .is_wysiwyg = "true";
defparam \stream_address[29] .power_up = "low";

dffeas \stream_address[30] (
	.clk(clk),
	.d(\Add0~121_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_30),
	.prn(vcc));
defparam \stream_address[30] .is_wysiwyg = "true";
defparam \stream_address[30] .power_up = "low";

dffeas \stream_address[31] (
	.clk(clk),
	.d(\Add0~125_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\stream_address~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(stream_address_31),
	.prn(vcc));
defparam \stream_address[31] .is_wysiwyg = "true";
defparam \stream_address[31] .power_up = "low";

dffeas \av_mif_addr[4] (
	.clk(clk),
	.d(\Add3~1_sumout ),
	.asdata(\mif_rec_addr[4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_4),
	.prn(vcc));
defparam \av_mif_addr[4] .is_wysiwyg = "true";
defparam \av_mif_addr[4] .power_up = "low";

dffeas \av_mif_addr[5] (
	.clk(clk),
	.d(\Add3~5_sumout ),
	.asdata(mif_rec_addr_5),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_5),
	.prn(vcc));
defparam \av_mif_addr[5] .is_wysiwyg = "true";
defparam \av_mif_addr[5] .power_up = "low";

dffeas \av_mif_addr[2] (
	.clk(clk),
	.d(\Add3~9_sumout ),
	.asdata(\mif_rec_addr[2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_2),
	.prn(vcc));
defparam \av_mif_addr[2] .is_wysiwyg = "true";
defparam \av_mif_addr[2] .power_up = "low";

dffeas \av_mif_addr[1] (
	.clk(clk),
	.d(\Add3~13_sumout ),
	.asdata(\mif_rec_addr[1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_1),
	.prn(vcc));
defparam \av_mif_addr[1] .is_wysiwyg = "true";
defparam \av_mif_addr[1] .power_up = "low";

dffeas \av_mif_addr[0] (
	.clk(clk),
	.d(\Add3~17_sumout ),
	.asdata(\mif_rec_addr[0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_0),
	.prn(vcc));
defparam \av_mif_addr[0] .is_wysiwyg = "true";
defparam \av_mif_addr[0] .power_up = "low";

dffeas \av_mif_addr[3] (
	.clk(clk),
	.d(\Add3~21_sumout ),
	.asdata(\mif_rec_addr[3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_3),
	.prn(vcc));
defparam \av_mif_addr[3] .is_wysiwyg = "true";
defparam \av_mif_addr[3] .power_up = "low";

dffeas \av_mif_addr[8] (
	.clk(clk),
	.d(\Add3~25_sumout ),
	.asdata(\mif_rec_addr[8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_8),
	.prn(vcc));
defparam \av_mif_addr[8] .is_wysiwyg = "true";
defparam \av_mif_addr[8] .power_up = "low";

dffeas \av_mif_addr[9] (
	.clk(clk),
	.d(\Add3~29_sumout ),
	.asdata(\mif_rec_addr[9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_9),
	.prn(vcc));
defparam \av_mif_addr[9] .is_wysiwyg = "true";
defparam \av_mif_addr[9] .power_up = "low";

dffeas \av_mif_addr[10] (
	.clk(clk),
	.d(\Add3~33_sumout ),
	.asdata(\mif_rec_addr[10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_10),
	.prn(vcc));
defparam \av_mif_addr[10] .is_wysiwyg = "true";
defparam \av_mif_addr[10] .power_up = "low";

dffeas \av_mif_addr[7] (
	.clk(clk),
	.d(\Add3~37_sumout ),
	.asdata(mif_rec_addr_7),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_7),
	.prn(vcc));
defparam \av_mif_addr[7] .is_wysiwyg = "true";
defparam \av_mif_addr[7] .power_up = "low";

dffeas \av_mif_addr[6] (
	.clk(clk),
	.d(\Add3~41_sumout ),
	.asdata(mif_rec_addr_6),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector2~1_combout ),
	.ena(\av_mif_addr[2]~3_combout ),
	.q(av_mif_addr_6),
	.prn(vcc));
defparam \av_mif_addr[6] .is_wysiwyg = "true";
defparam \av_mif_addr[6] .power_up = "low";

dffeas stream_read(
	.clk(clk),
	.d(\stream_read~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stream_read1),
	.prn(vcc));
defparam stream_read.is_wysiwyg = "true";
defparam stream_read.power_up = "low";

dffeas av_ctrl_req(
	.clk(clk),
	.d(\av_ctrl_req~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_ctrl_req1),
	.prn(vcc));
defparam av_ctrl_req.is_wysiwyg = "true";
defparam av_ctrl_req.power_up = "low";

dffeas pll_go(
	.clk(clk),
	.d(\pll_go~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pll_go1),
	.prn(vcc));
defparam pll_go.is_wysiwyg = "true";
defparam pll_go.power_up = "low";

dffeas av_addr_burst(
	.clk(clk),
	.d(\Equal0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_addr_burst1),
	.prn(vcc));
defparam av_addr_burst.is_wysiwyg = "true";
defparam av_addr_burst.power_up = "low";

dffeas av_opcode_err(
	.clk(clk),
	.d(\av_opcode_err~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_opcode_err1),
	.prn(vcc));
defparam av_opcode_err.is_wysiwyg = "true";
defparam av_opcode_err.power_up = "low";

dffeas av_done(
	.clk(clk),
	.d(\av_done~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_done1),
	.prn(vcc));
defparam av_done.is_wysiwyg = "true";
defparam av_done.power_up = "low";

dffeas pll_type(
	.clk(clk),
	.d(\rec_is_cgb~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pll_type1),
	.prn(vcc));
defparam pll_type.is_wysiwyg = "true";
defparam pll_type.power_up = "low";

dffeas \mif_rec_data[1] (
	.clk(clk),
	.d(stream_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_1),
	.prn(vcc));
defparam \mif_rec_data[1] .is_wysiwyg = "true";
defparam \mif_rec_data[1] .power_up = "low";

dffeas \mif_rec_addr[7] (
	.clk(clk),
	.d(stream_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(mif_rec_addr_7),
	.prn(vcc));
defparam \mif_rec_addr[7] .is_wysiwyg = "true";
defparam \mif_rec_addr[7] .power_up = "low";

dffeas \mif_rec_addr[5] (
	.clk(clk),
	.d(stream_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(mif_rec_addr_5),
	.prn(vcc));
defparam \mif_rec_addr[5] .is_wysiwyg = "true";
defparam \mif_rec_addr[5] .power_up = "low";

dffeas \mif_rec_addr[6] (
	.clk(clk),
	.d(stream_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(mif_rec_addr_6),
	.prn(vcc));
defparam \mif_rec_addr[6] .is_wysiwyg = "true";
defparam \mif_rec_addr[6] .power_up = "low";

dffeas \mif_rec_data[2] (
	.clk(clk),
	.d(stream_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_2),
	.prn(vcc));
defparam \mif_rec_data[2] .is_wysiwyg = "true";
defparam \mif_rec_data[2] .power_up = "low";

dffeas \mif_rec_data[0] (
	.clk(clk),
	.d(stream_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_0),
	.prn(vcc));
defparam \mif_rec_data[0] .is_wysiwyg = "true";
defparam \mif_rec_data[0] .power_up = "low";

dffeas \mif_rec_data[3] (
	.clk(clk),
	.d(stream_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_3),
	.prn(vcc));
defparam \mif_rec_data[3] .is_wysiwyg = "true";
defparam \mif_rec_data[3] .power_up = "low";

dffeas av_mif_type_valid(
	.clk(clk),
	.d(\rec_is_type~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_mif_type_valid1),
	.prn(vcc));
defparam av_mif_type_valid.is_wysiwyg = "true";
defparam av_mif_type_valid.power_up = "low";

dffeas \av_mif_type[1] (
	.clk(clk),
	.d(\av_mif_type~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_mif_type_1),
	.prn(vcc));
defparam \av_mif_type[1] .is_wysiwyg = "true";
defparam \av_mif_type[1] .power_up = "low";

dffeas \av_mif_type[0] (
	.clk(clk),
	.d(\av_mif_type~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_mif_type_0),
	.prn(vcc));
defparam \av_mif_type[0] .is_wysiwyg = "true";
defparam \av_mif_type[0] .power_up = "low";

dffeas \mif_rec_data[4] (
	.clk(clk),
	.d(stream_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_4),
	.prn(vcc));
defparam \mif_rec_data[4] .is_wysiwyg = "true";
defparam \mif_rec_data[4] .power_up = "low";

dffeas \mif_rec_data[5] (
	.clk(clk),
	.d(stream_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_5),
	.prn(vcc));
defparam \mif_rec_data[5] .is_wysiwyg = "true";
defparam \mif_rec_data[5] .power_up = "low";

dffeas \mif_rec_data[6] (
	.clk(clk),
	.d(stream_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_6),
	.prn(vcc));
defparam \mif_rec_data[6] .is_wysiwyg = "true";
defparam \mif_rec_data[6] .power_up = "low";

dffeas \mif_rec_data[7] (
	.clk(clk),
	.d(stream_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_7),
	.prn(vcc));
defparam \mif_rec_data[7] .is_wysiwyg = "true";
defparam \mif_rec_data[7] .power_up = "low";

dffeas \mif_rec_data[8] (
	.clk(clk),
	.d(stream_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_8),
	.prn(vcc));
defparam \mif_rec_data[8] .is_wysiwyg = "true";
defparam \mif_rec_data[8] .power_up = "low";

dffeas \mif_rec_data[9] (
	.clk(clk),
	.d(stream_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_9),
	.prn(vcc));
defparam \mif_rec_data[9] .is_wysiwyg = "true";
defparam \mif_rec_data[9] .power_up = "low";

dffeas \mif_rec_data[10] (
	.clk(clk),
	.d(stream_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_10),
	.prn(vcc));
defparam \mif_rec_data[10] .is_wysiwyg = "true";
defparam \mif_rec_data[10] .power_up = "low";

dffeas \mif_rec_data[11] (
	.clk(clk),
	.d(stream_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_11),
	.prn(vcc));
defparam \mif_rec_data[11] .is_wysiwyg = "true";
defparam \mif_rec_data[11] .power_up = "low";

dffeas \mif_rec_data[12] (
	.clk(clk),
	.d(stream_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_12),
	.prn(vcc));
defparam \mif_rec_data[12] .is_wysiwyg = "true";
defparam \mif_rec_data[12] .power_up = "low";

dffeas \mif_rec_data[13] (
	.clk(clk),
	.d(stream_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_13),
	.prn(vcc));
defparam \mif_rec_data[13] .is_wysiwyg = "true";
defparam \mif_rec_data[13] .power_up = "low";

dffeas \mif_rec_data[14] (
	.clk(clk),
	.d(stream_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_14),
	.prn(vcc));
defparam \mif_rec_data[14] .is_wysiwyg = "true";
defparam \mif_rec_data[14] .power_up = "low";

dffeas \mif_rec_data[15] (
	.clk(clk),
	.d(stream_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_rec_data~0_combout ),
	.q(mif_rec_data_15),
	.prn(vcc));
defparam \mif_rec_data[15] .is_wysiwyg = "true";
defparam \mif_rec_data[15] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[0]~q ),
	.datae(gnd),
	.dataf(!mif_addr_mode),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~1 .shared_arith = "off";

dffeas \av_state.AV_DEC_HDR (
	.clk(clk),
	.d(\av_next_state.AV_DEC_HDR~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_state.AV_DEC_HDR~q ),
	.prn(vcc));
defparam \av_state.AV_DEC_HDR .is_wysiwyg = "true";
defparam \av_state.AV_DEC_HDR .power_up = "low";

dffeas \mif_rec_len[0] (
	.clk(clk),
	.d(stream_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_len[0]~q ),
	.prn(vcc));
defparam \mif_rec_len[0] .is_wysiwyg = "true";
defparam \mif_rec_len[0] .power_up = "low";

dffeas \mif_rec_len[4] (
	.clk(clk),
	.d(stream_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_len[4]~q ),
	.prn(vcc));
defparam \mif_rec_len[4] .is_wysiwyg = "true";
defparam \mif_rec_len[4] .power_up = "low";

dffeas \mif_rec_len[3] (
	.clk(clk),
	.d(stream_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_len[3]~q ),
	.prn(vcc));
defparam \mif_rec_len[3] .is_wysiwyg = "true";
defparam \mif_rec_len[3] .power_up = "low";

dffeas \mif_rec_len[2] (
	.clk(clk),
	.d(stream_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_len[2]~q ),
	.prn(vcc));
defparam \mif_rec_len[2] .is_wysiwyg = "true";
defparam \mif_rec_len[2] .power_up = "low";

dffeas \mif_rec_len[1] (
	.clk(clk),
	.d(stream_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_len[1]~q ),
	.prn(vcc));
defparam \mif_rec_len[1] .is_wysiwyg = "true";
defparam \mif_rec_len[1] .power_up = "low";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!\mif_rec_len[4]~q ),
	.datab(!\mif_rec_len[3]~q ),
	.datac(!\mif_rec_len[2]~q ),
	.datad(!\mif_rec_len[1]~q ),
	.datae(!\mif_rec_len[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h8000000080000000;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_len_cnt[1]~7 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\mif_len_cnt[1]~q ),
	.datac(!\av_state.AV_DEC_HDR~q ),
	.datad(!\mif_rec_len[1]~q ),
	.datae(!\Equal2~0_combout ),
	.dataf(!\mif_len_cnt[4]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[1]~7 .extended_lut = "off";
defparam \mif_len_cnt[1]~7 .lut_mask = 64'h909F999F33333333;
defparam \mif_len_cnt[1]~7 .shared_arith = "off";

dffeas \mif_len_cnt[1] (
	.clk(clk),
	.d(\mif_len_cnt[1]~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mif_len_cnt[1]~q ),
	.prn(vcc));
defparam \mif_len_cnt[1] .is_wysiwyg = "true";
defparam \mif_len_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!\av_state.AV_DEC_HDR~q ),
	.datab(!\Equal2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h4444444444444444;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \mif_len_cnt[2]~5 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\mif_len_cnt[2]~q ),
	.datac(!\mif_len_cnt[1]~q ),
	.datad(!\Selector2~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[2]~5 .extended_lut = "off";
defparam \mif_len_cnt[2]~5 .lut_mask = 64'h9300930093009300;
defparam \mif_len_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \mif_len_cnt[2]~6 (
	.dataa(!\mif_len_cnt[2]~q ),
	.datab(!\av_state.AV_DEC_HDR~q ),
	.datac(!\mif_rec_len[2]~q ),
	.datad(!\mif_len_cnt[4]~0_combout ),
	.datae(!\mif_len_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[2]~6 .extended_lut = "off";
defparam \mif_len_cnt[2]~6 .lut_mask = 64'h0355FF550355FF55;
defparam \mif_len_cnt[2]~6 .shared_arith = "off";

dffeas \mif_len_cnt[2] (
	.clk(clk),
	.d(\mif_len_cnt[2]~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mif_len_cnt[2]~q ),
	.prn(vcc));
defparam \mif_len_cnt[2] .is_wysiwyg = "true";
defparam \mif_len_cnt[2] .power_up = "low";

cyclonev_lcell_comb \mif_len_cnt[3]~3 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\mif_len_cnt[3]~q ),
	.datac(!\mif_len_cnt[2]~q ),
	.datad(!\mif_len_cnt[1]~q ),
	.datae(!\Selector2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[3]~3 .extended_lut = "off";
defparam \mif_len_cnt[3]~3 .lut_mask = 64'h9333000093330000;
defparam \mif_len_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \mif_len_cnt[3]~4 (
	.dataa(!\mif_len_cnt[3]~q ),
	.datab(!\av_state.AV_DEC_HDR~q ),
	.datac(!\mif_rec_len[3]~q ),
	.datad(!\mif_len_cnt[4]~0_combout ),
	.datae(!\mif_len_cnt[3]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[3]~4 .extended_lut = "off";
defparam \mif_len_cnt[3]~4 .lut_mask = 64'h0355FF550355FF55;
defparam \mif_len_cnt[3]~4 .shared_arith = "off";

dffeas \mif_len_cnt[3] (
	.clk(clk),
	.d(\mif_len_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mif_len_cnt[3]~q ),
	.prn(vcc));
defparam \mif_len_cnt[3] .is_wysiwyg = "true";
defparam \mif_len_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\mif_len_cnt[3]~q ),
	.datac(!\mif_len_cnt[2]~q ),
	.datad(!\mif_len_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h8000800080008000;
defparam \Add2~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_len_cnt[4]~2 (
	.dataa(!\mif_len_cnt[4]~q ),
	.datab(!\av_state.AV_DEC_HDR~q ),
	.datac(!\mif_rec_len[4]~q ),
	.datad(!\Equal2~0_combout ),
	.datae(!\mif_len_cnt[4]~0_combout ),
	.dataf(!\Add2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[4]~2 .extended_lut = "off";
defparam \mif_len_cnt[4]~2 .lut_mask = 64'h475755558BAB5555;
defparam \mif_len_cnt[4]~2 .shared_arith = "off";

dffeas \mif_len_cnt[4] (
	.clk(clk),
	.d(\mif_len_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mif_len_cnt[4]~q ),
	.prn(vcc));
defparam \mif_len_cnt[4] .is_wysiwyg = "true";
defparam \mif_len_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\mif_len_cnt[4]~q ),
	.datab(!\mif_len_cnt[3]~q ),
	.datac(!\mif_len_cnt[2]~q ),
	.datad(!\mif_len_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal0~0 .shared_arith = "off";

dffeas \mif_rec_addr[1] (
	.clk(clk),
	.d(stream_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[1]~q ),
	.prn(vcc));
defparam \mif_rec_addr[1] .is_wysiwyg = "true";
defparam \mif_rec_addr[1] .power_up = "low";

dffeas \mif_rec_addr[0] (
	.clk(clk),
	.d(stream_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[0]~q ),
	.prn(vcc));
defparam \mif_rec_addr[0] .is_wysiwyg = "true";
defparam \mif_rec_addr[0] .power_up = "low";

dffeas \mif_rec_addr[4] (
	.clk(clk),
	.d(stream_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[4]~q ),
	.prn(vcc));
defparam \mif_rec_addr[4] .is_wysiwyg = "true";
defparam \mif_rec_addr[4] .power_up = "low";

dffeas \mif_rec_addr[3] (
	.clk(clk),
	.d(stream_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[3]~q ),
	.prn(vcc));
defparam \mif_rec_addr[3] .is_wysiwyg = "true";
defparam \mif_rec_addr[3] .power_up = "low";

dffeas \mif_rec_addr[2] (
	.clk(clk),
	.d(stream_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[2]~q ),
	.prn(vcc));
defparam \mif_rec_addr[2] .is_wysiwyg = "true";
defparam \mif_rec_addr[2] .power_up = "low";

cyclonev_lcell_comb \rec_is_eom~0 (
	.dataa(!\mif_rec_addr[4]~q ),
	.datab(!\mif_rec_addr[3]~q ),
	.datac(!\mif_rec_addr[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rec_is_eom~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rec_is_eom~0 .extended_lut = "off";
defparam \rec_is_eom~0 .lut_mask = 64'h0101010101010101;
defparam \rec_is_eom~0 .shared_arith = "off";

cyclonev_lcell_comb \rec_is_eom~1 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\av_state.AV_IDLE~q ),
	.datac(!\mif_rec_addr[1]~q ),
	.datad(!\mif_rec_addr[0]~q ),
	.datae(!\rec_is_eom~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rec_is_eom~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rec_is_eom~1 .extended_lut = "off";
defparam \rec_is_eom~1 .lut_mask = 64'h0000000100000001;
defparam \rec_is_eom~1 .shared_arith = "off";

cyclonev_lcell_comb \invalid_rec~0 (
	.dataa(!\mif_rec_addr[4]~q ),
	.datab(!\mif_rec_addr[3]~q ),
	.datac(!\mif_rec_addr[2]~q ),
	.datad(!\mif_rec_addr[1]~q ),
	.datae(!\mif_rec_addr[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\invalid_rec~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \invalid_rec~0 .extended_lut = "off";
defparam \invalid_rec~0 .lut_mask = 64'h0800008008000080;
defparam \invalid_rec~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_strm_active~0 (
	.dataa(!\av_next_state.AV_DEC_HDR~0_combout ),
	.datab(!\mif_strm_active~q ),
	.datac(!\Selector0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_strm_active~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_strm_active~0 .extended_lut = "off";
defparam \mif_strm_active~0 .lut_mask = 64'h5757575757575757;
defparam \mif_strm_active~0 .shared_arith = "off";

dffeas mif_strm_active(
	.clk(clk),
	.d(\mif_strm_active~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mif_strm_active~q ),
	.prn(vcc));
defparam mif_strm_active.is_wysiwyg = "true";
defparam mif_strm_active.power_up = "low";

cyclonev_lcell_comb \invalid_rec~1 (
	.dataa(!\mif_rec_addr[4]~q ),
	.datab(!\mif_rec_addr[3]~q ),
	.datac(!\mif_rec_addr[2]~q ),
	.datad(!\mif_rec_addr[1]~q ),
	.datae(!\mif_rec_addr[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\invalid_rec~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \invalid_rec~1 .extended_lut = "off";
defparam \invalid_rec~1 .lut_mask = 64'h0880808108808081;
defparam \invalid_rec~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~1 (
	.dataa(!\av_state.AV_DEC_HDR~q ),
	.datab(!\Equal2~0_combout ),
	.datac(!\invalid_rec~0_combout ),
	.datad(!\mif_strm_active~q ),
	.datae(!\invalid_rec~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'h0010000000100000;
defparam \Selector4~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~2 (
	.dataa(!mif_err_reg_4),
	.datab(!mif_err_reg_1),
	.datac(!mif_err_reg_0),
	.datad(!\Selector4~0_combout ),
	.datae(!\Selector4~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~2 .extended_lut = "off";
defparam \Selector4~2 .lut_mask = 64'h007FFFFF007FFFFF;
defparam \Selector4~2 .shared_arith = "off";

dffeas \av_state.AV_REC_ERR (
	.clk(clk),
	.d(\Selector4~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_state.AV_REC_ERR~q ),
	.prn(vcc));
defparam \av_state.AV_REC_ERR .is_wysiwyg = "true";
defparam \av_state.AV_REC_ERR .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\av_state.AV_DEC_HDR~q ),
	.datab(!ctrl_av_go),
	.datac(!\av_state.AV_IDLE~q ),
	.datad(!\rec_is_eom~1_combout ),
	.datae(!\av_state.AV_REC_ERR~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h3F2A00003F2A0000;
defparam \Selector0~0 .shared_arith = "off";

dffeas \av_state.AV_IDLE (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_state.AV_IDLE~q ),
	.prn(vcc));
defparam \av_state.AV_IDLE .is_wysiwyg = "true";
defparam \av_state.AV_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector3~3 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!ctrl_op_done),
	.datad(!\Selector3~2_combout ),
	.datae(!\mif_rec_data~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~3 .extended_lut = "off";
defparam \Selector3~3 .lut_mask = 64'hFF0F8808FF0F8808;
defparam \Selector3~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~4 (
	.dataa(!\av_state.AV_DEC_HDR~q ),
	.datab(!\Equal2~0_combout ),
	.datac(!\av_state.AV_IDLE~q ),
	.datad(!\invalid_rec~0_combout ),
	.datae(!\Selector3~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~4 .extended_lut = "off";
defparam \Selector3~4 .lut_mask = 64'hFFFF0001FFFF0001;
defparam \Selector3~4 .shared_arith = "off";

dffeas \av_state.AV_WF_DONE (
	.clk(clk),
	.d(\Selector3~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_state.AV_WF_DONE~q ),
	.prn(vcc));
defparam \av_state.AV_WF_DONE .is_wysiwyg = "true";
defparam \av_state.AV_WF_DONE .power_up = "low";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!pll_mif_busy),
	.datab(!\pll_active_dly~q ),
	.datac(!\av_state.AV_WF_DONE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h0202020202020202;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \pll_active~0 (
	.dataa(!\av_state.AV_DEC_HDR~q ),
	.datab(!\Equal2~0_combout ),
	.datac(!\av_state.AV_IDLE~q ),
	.datad(!\Selector1~2_combout ),
	.datae(!\invalid_rec~0_combout ),
	.dataf(!\pll_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_active~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_active~0 .extended_lut = "off";
defparam \pll_active~0 .lut_mask = 64'h00000101FF00FF01;
defparam \pll_active~0 .shared_arith = "off";

dffeas pll_active(
	.clk(clk),
	.d(\pll_active~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_active~q ),
	.prn(vcc));
defparam pll_active.is_wysiwyg = "true";
defparam pll_active.power_up = "low";

dffeas pll_active_dly(
	.clk(clk),
	.d(\pll_active~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_active_dly~q ),
	.prn(vcc));
defparam pll_active_dly.is_wysiwyg = "true";
defparam pll_active_dly.power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!pll_mif_busy),
	.datab(!\pll_active_dly~q ),
	.datac(!\av_state.AV_WF_DONE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h0D0D0D0D0D0D0D0D;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~2 (
	.dataa(!mif_err_reg_4),
	.datab(!mif_err_reg_1),
	.datac(!mif_err_reg_0),
	.datad(!\Selector4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~2 .extended_lut = "off";
defparam \Selector3~2 .lut_mask = 64'h0080008000800080;
defparam \Selector3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!stream_read1),
	.datab(!reconfig_mif_waitrequest),
	.datac(!\mif_len_cnt[0]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\av_state.AV_RD_DATA~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'h00000BBB00000BBB;
defparam \Selector2~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~3 (
	.dataa(!\Selector2~1_combout ),
	.datab(!ctrl_op_done),
	.datac(!\Selector3~2_combout ),
	.datad(!\Selector2~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~3 .extended_lut = "off";
defparam \Selector2~3 .lut_mask = 64'h57FF57FF57FF57FF;
defparam \Selector2~3 .shared_arith = "off";

dffeas \av_state.AV_RD_DATA (
	.clk(clk),
	.d(\Selector2~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_state.AV_RD_DATA~q ),
	.prn(vcc));
defparam \av_state.AV_RD_DATA .is_wysiwyg = "true";
defparam \av_state.AV_RD_DATA .power_up = "low";

cyclonev_lcell_comb \mif_rec_data~0 (
	.dataa(!stream_read1),
	.datab(!reconfig_mif_waitrequest),
	.datac(!\av_state.AV_RD_DATA~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_rec_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_rec_data~0 .extended_lut = "off";
defparam \mif_rec_data~0 .lut_mask = 64'h0404040404040404;
defparam \mif_rec_data~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_len_cnt[4]~0 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!\Selector2~1_combout ),
	.datad(!\mif_rec_data~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[4]~0 .extended_lut = "off";
defparam \mif_len_cnt[4]~0 .lut_mask = 64'hF080F080F080F080;
defparam \mif_len_cnt[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_len_cnt[0]~1 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\av_state.AV_DEC_HDR~q ),
	.datac(!\mif_rec_len[0]~q ),
	.datad(!\Equal2~0_combout ),
	.datae(!\mif_len_cnt[4]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_len_cnt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_len_cnt[0]~1 .extended_lut = "off";
defparam \mif_len_cnt[0]~1 .lut_mask = 64'h8BAB55558BAB5555;
defparam \mif_len_cnt[0]~1 .shared_arith = "off";

dffeas \mif_len_cnt[0] (
	.clk(clk),
	.d(\mif_len_cnt[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mif_len_cnt[0]~q ),
	.prn(vcc));
defparam \mif_len_cnt[0] .is_wysiwyg = "true";
defparam \mif_len_cnt[0] .power_up = "low";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!\mif_rec_addr[4]~q ),
	.datab(!\mif_rec_addr[3]~q ),
	.datac(!\mif_rec_addr[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h8080808080808080;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \rec_is_som~0 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\av_state.AV_IDLE~q ),
	.datac(!\mif_rec_addr[1]~q ),
	.datad(!\mif_rec_addr[0]~q ),
	.datae(!\Equal6~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rec_is_som~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rec_is_som~0 .extended_lut = "off";
defparam \rec_is_som~0 .lut_mask = 64'h0000001000000010;
defparam \rec_is_som~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\av_state.AV_IDLE~q ),
	.datac(!\invalid_rec~0_combout ),
	.datad(!\mif_strm_active~q ),
	.datae(!\invalid_rec~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h5400541054005410;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~4 (
	.dataa(!\av_state.AV_DEC_HDR~q ),
	.datab(!\rec_is_eom~1_combout ),
	.datac(!\rec_is_som~0_combout ),
	.datad(!\Selector1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~4 .extended_lut = "off";
defparam \Selector1~4 .lut_mask = 64'h0444044404440444;
defparam \Selector1~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~5 (
	.dataa(!stream_read1),
	.datab(!reconfig_mif_waitrequest),
	.datac(!\av_state.AV_RD_HDR~q ),
	.datad(!ctrl_av_go),
	.datae(!\av_state.AV_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~5 .extended_lut = "off";
defparam \Selector1~5 .lut_mask = 64'hF400F4F4F400F4F4;
defparam \Selector1~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~7 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!\av_state.AV_RD_DATA~q ),
	.datad(!\Selector1~2_combout ),
	.datae(!\Selector1~4_combout ),
	.dataf(!\Selector1~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~7 .extended_lut = "off";
defparam \Selector1~7 .lut_mask = 64'hFFFFFFFF08FFFFFF;
defparam \Selector1~7 .shared_arith = "off";

dffeas \av_state.AV_RD_HDR (
	.clk(clk),
	.d(\Selector1~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_state.AV_RD_HDR~q ),
	.prn(vcc));
defparam \av_state.AV_RD_HDR .is_wysiwyg = "true";
defparam \av_state.AV_RD_HDR .power_up = "low";

cyclonev_lcell_comb \av_next_state.AV_DEC_HDR~0 (
	.dataa(!stream_read1),
	.datab(!reconfig_mif_waitrequest),
	.datac(!\av_state.AV_RD_HDR~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_next_state.AV_DEC_HDR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_next_state.AV_DEC_HDR~0 .extended_lut = "off";
defparam \av_next_state.AV_DEC_HDR~0 .lut_mask = 64'h0404040404040404;
defparam \av_next_state.AV_DEC_HDR~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_next_offset~0 (
	.dataa(!\av_next_state.AV_DEC_HDR~0_combout ),
	.datab(!\mif_len_cnt[0]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\mif_rec_data~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_next_offset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_next_offset~0 .extended_lut = "off";
defparam \mif_next_offset~0 .lut_mask = 64'hAA80AA80AA80AA80;
defparam \mif_next_offset~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_next_offset[28]~1 (
	.dataa(!\Selector0~0_combout ),
	.datab(!\mif_next_offset~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_next_offset[28]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_next_offset[28]~1 .extended_lut = "off";
defparam \mif_next_offset[28]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \mif_next_offset[28]~1 .shared_arith = "off";

dffeas \mif_next_offset[0] (
	.clk(clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[0]~q ),
	.prn(vcc));
defparam \mif_next_offset[0] .is_wysiwyg = "true";
defparam \mif_next_offset[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[0]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~6 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!\av_state.AV_RD_DATA~q ),
	.datad(!\Selector1~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~6 .extended_lut = "off";
defparam \Selector1~6 .lut_mask = 64'h00F700F700F700F7;
defparam \Selector1~6 .shared_arith = "off";

cyclonev_lcell_comb \stream_address~0 (
	.dataa(!\av_next_state.AV_DEC_HDR~0_combout ),
	.datab(!\Selector1~2_combout ),
	.datac(!\Selector2~3_combout ),
	.datad(!\Selector1~4_combout ),
	.datae(!\Selector1~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stream_address~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stream_address~0 .extended_lut = "off";
defparam \stream_address~0 .lut_mask = 64'h0000800000008000;
defparam \stream_address~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[1]~q ),
	.datae(gnd),
	.dataf(!mif_addr_mode),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000FF000000FF;
defparam \Add1~5 .shared_arith = "off";

dffeas \mif_next_offset[1] (
	.clk(clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[1]~q ),
	.prn(vcc));
defparam \mif_next_offset[1] .is_wysiwyg = "true";
defparam \mif_next_offset[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[1]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_1),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

dffeas \mif_next_offset[2] (
	.clk(clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[2]~q ),
	.prn(vcc));
defparam \mif_next_offset[2] .is_wysiwyg = "true";
defparam \mif_next_offset[2] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[2]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_2),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

dffeas \mif_next_offset[3] (
	.clk(clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[3]~q ),
	.prn(vcc));
defparam \mif_next_offset[3] .is_wysiwyg = "true";
defparam \mif_next_offset[3] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[3]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_3),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

dffeas \mif_next_offset[4] (
	.clk(clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[4]~q ),
	.prn(vcc));
defparam \mif_next_offset[4] .is_wysiwyg = "true";
defparam \mif_next_offset[4] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[4]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_4),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

dffeas \mif_next_offset[5] (
	.clk(clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[5]~q ),
	.prn(vcc));
defparam \mif_next_offset[5] .is_wysiwyg = "true";
defparam \mif_next_offset[5] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[5]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_5),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~25 .shared_arith = "off";

dffeas \mif_next_offset[6] (
	.clk(clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[6]~q ),
	.prn(vcc));
defparam \mif_next_offset[6] .is_wysiwyg = "true";
defparam \mif_next_offset[6] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[6]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_6),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~29 .shared_arith = "off";

dffeas \mif_next_offset[7] (
	.clk(clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[7]~q ),
	.prn(vcc));
defparam \mif_next_offset[7] .is_wysiwyg = "true";
defparam \mif_next_offset[7] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[7]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_7),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~33 .shared_arith = "off";

dffeas \mif_next_offset[8] (
	.clk(clk),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[8]~q ),
	.prn(vcc));
defparam \mif_next_offset[8] .is_wysiwyg = "true";
defparam \mif_next_offset[8] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[8]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_8),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout());
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~37 .shared_arith = "off";

dffeas \mif_next_offset[9] (
	.clk(clk),
	.d(\Add1~37_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[9]~q ),
	.prn(vcc));
defparam \mif_next_offset[9] .is_wysiwyg = "true";
defparam \mif_next_offset[9] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[9]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_9),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(\Add1~42 ),
	.shareout());
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~41 .shared_arith = "off";

dffeas \mif_next_offset[10] (
	.clk(clk),
	.d(\Add1~41_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[10]~q ),
	.prn(vcc));
defparam \mif_next_offset[10] .is_wysiwyg = "true";
defparam \mif_next_offset[10] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[10]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_10),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~45_sumout ),
	.cout(\Add1~46 ),
	.shareout());
defparam \Add1~45 .extended_lut = "off";
defparam \Add1~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~45 .shared_arith = "off";

dffeas \mif_next_offset[11] (
	.clk(clk),
	.d(\Add1~45_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[11]~q ),
	.prn(vcc));
defparam \mif_next_offset[11] .is_wysiwyg = "true";
defparam \mif_next_offset[11] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[11]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_11),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~49_sumout ),
	.cout(\Add1~50 ),
	.shareout());
defparam \Add1~49 .extended_lut = "off";
defparam \Add1~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~49 .shared_arith = "off";

dffeas \mif_next_offset[12] (
	.clk(clk),
	.d(\Add1~49_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[12]~q ),
	.prn(vcc));
defparam \mif_next_offset[12] .is_wysiwyg = "true";
defparam \mif_next_offset[12] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[12]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_12),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \Add1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~53_sumout ),
	.cout(\Add1~54 ),
	.shareout());
defparam \Add1~53 .extended_lut = "off";
defparam \Add1~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~53 .shared_arith = "off";

dffeas \mif_next_offset[13] (
	.clk(clk),
	.d(\Add1~53_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[13]~q ),
	.prn(vcc));
defparam \mif_next_offset[13] .is_wysiwyg = "true";
defparam \mif_next_offset[13] .power_up = "low";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[13]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_13),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \Add1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~57_sumout ),
	.cout(\Add1~58 ),
	.shareout());
defparam \Add1~57 .extended_lut = "off";
defparam \Add1~57 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~57 .shared_arith = "off";

dffeas \mif_next_offset[14] (
	.clk(clk),
	.d(\Add1~57_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[14]~q ),
	.prn(vcc));
defparam \mif_next_offset[14] .is_wysiwyg = "true";
defparam \mif_next_offset[14] .power_up = "low";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[14]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_14),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \Add1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~61_sumout ),
	.cout(\Add1~62 ),
	.shareout());
defparam \Add1~61 .extended_lut = "off";
defparam \Add1~61 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~61 .shared_arith = "off";

dffeas \mif_next_offset[15] (
	.clk(clk),
	.d(\Add1~61_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[15]~q ),
	.prn(vcc));
defparam \mif_next_offset[15] .is_wysiwyg = "true";
defparam \mif_next_offset[15] .power_up = "low";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[15]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_15),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \Add1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~65_sumout ),
	.cout(\Add1~66 ),
	.shareout());
defparam \Add1~65 .extended_lut = "off";
defparam \Add1~65 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~65 .shared_arith = "off";

dffeas \mif_next_offset[16] (
	.clk(clk),
	.d(\Add1~65_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[16]~q ),
	.prn(vcc));
defparam \mif_next_offset[16] .is_wysiwyg = "true";
defparam \mif_next_offset[16] .power_up = "low";

cyclonev_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[16]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_16),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

cyclonev_lcell_comb \Add1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~69_sumout ),
	.cout(\Add1~70 ),
	.shareout());
defparam \Add1~69 .extended_lut = "off";
defparam \Add1~69 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~69 .shared_arith = "off";

dffeas \mif_next_offset[17] (
	.clk(clk),
	.d(\Add1~69_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[17]~q ),
	.prn(vcc));
defparam \mif_next_offset[17] .is_wysiwyg = "true";
defparam \mif_next_offset[17] .power_up = "low";

cyclonev_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[17]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_17),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

cyclonev_lcell_comb \Add1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~73_sumout ),
	.cout(\Add1~74 ),
	.shareout());
defparam \Add1~73 .extended_lut = "off";
defparam \Add1~73 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~73 .shared_arith = "off";

dffeas \mif_next_offset[18] (
	.clk(clk),
	.d(\Add1~73_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[18]~q ),
	.prn(vcc));
defparam \mif_next_offset[18] .is_wysiwyg = "true";
defparam \mif_next_offset[18] .power_up = "low";

cyclonev_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[18]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_18),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

cyclonev_lcell_comb \Add1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~77_sumout ),
	.cout(\Add1~78 ),
	.shareout());
defparam \Add1~77 .extended_lut = "off";
defparam \Add1~77 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~77 .shared_arith = "off";

dffeas \mif_next_offset[19] (
	.clk(clk),
	.d(\Add1~77_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[19]~q ),
	.prn(vcc));
defparam \mif_next_offset[19] .is_wysiwyg = "true";
defparam \mif_next_offset[19] .power_up = "low";

cyclonev_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[19]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_19),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

cyclonev_lcell_comb \Add1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~81_sumout ),
	.cout(\Add1~82 ),
	.shareout());
defparam \Add1~81 .extended_lut = "off";
defparam \Add1~81 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~81 .shared_arith = "off";

dffeas \mif_next_offset[20] (
	.clk(clk),
	.d(\Add1~81_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[20]~q ),
	.prn(vcc));
defparam \mif_next_offset[20] .is_wysiwyg = "true";
defparam \mif_next_offset[20] .power_up = "low";

cyclonev_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[20]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_20),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

cyclonev_lcell_comb \Add1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~85_sumout ),
	.cout(\Add1~86 ),
	.shareout());
defparam \Add1~85 .extended_lut = "off";
defparam \Add1~85 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~85 .shared_arith = "off";

dffeas \mif_next_offset[21] (
	.clk(clk),
	.d(\Add1~85_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[21]~q ),
	.prn(vcc));
defparam \mif_next_offset[21] .is_wysiwyg = "true";
defparam \mif_next_offset[21] .power_up = "low";

cyclonev_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[21]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_21),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

cyclonev_lcell_comb \Add1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~89_sumout ),
	.cout(\Add1~90 ),
	.shareout());
defparam \Add1~89 .extended_lut = "off";
defparam \Add1~89 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~89 .shared_arith = "off";

dffeas \mif_next_offset[22] (
	.clk(clk),
	.d(\Add1~89_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[22]~q ),
	.prn(vcc));
defparam \mif_next_offset[22] .is_wysiwyg = "true";
defparam \mif_next_offset[22] .power_up = "low";

cyclonev_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[22]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_22),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

cyclonev_lcell_comb \Add1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~93_sumout ),
	.cout(\Add1~94 ),
	.shareout());
defparam \Add1~93 .extended_lut = "off";
defparam \Add1~93 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~93 .shared_arith = "off";

dffeas \mif_next_offset[23] (
	.clk(clk),
	.d(\Add1~93_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[23]~q ),
	.prn(vcc));
defparam \mif_next_offset[23] .is_wysiwyg = "true";
defparam \mif_next_offset[23] .power_up = "low";

cyclonev_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[23]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_23),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

cyclonev_lcell_comb \Add1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~97_sumout ),
	.cout(\Add1~98 ),
	.shareout());
defparam \Add1~97 .extended_lut = "off";
defparam \Add1~97 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~97 .shared_arith = "off";

dffeas \mif_next_offset[24] (
	.clk(clk),
	.d(\Add1~97_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[24]~q ),
	.prn(vcc));
defparam \mif_next_offset[24] .is_wysiwyg = "true";
defparam \mif_next_offset[24] .power_up = "low";

cyclonev_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[24]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_24),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

cyclonev_lcell_comb \Add1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~101_sumout ),
	.cout(\Add1~102 ),
	.shareout());
defparam \Add1~101 .extended_lut = "off";
defparam \Add1~101 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~101 .shared_arith = "off";

dffeas \mif_next_offset[25] (
	.clk(clk),
	.d(\Add1~101_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[25]~q ),
	.prn(vcc));
defparam \mif_next_offset[25] .is_wysiwyg = "true";
defparam \mif_next_offset[25] .power_up = "low";

cyclonev_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[25]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_25),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

cyclonev_lcell_comb \Add1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~105_sumout ),
	.cout(\Add1~106 ),
	.shareout());
defparam \Add1~105 .extended_lut = "off";
defparam \Add1~105 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~105 .shared_arith = "off";

dffeas \mif_next_offset[26] (
	.clk(clk),
	.d(\Add1~105_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[26]~q ),
	.prn(vcc));
defparam \mif_next_offset[26] .is_wysiwyg = "true";
defparam \mif_next_offset[26] .power_up = "low";

cyclonev_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[26]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_26),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

cyclonev_lcell_comb \Add1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~109_sumout ),
	.cout(\Add1~110 ),
	.shareout());
defparam \Add1~109 .extended_lut = "off";
defparam \Add1~109 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~109 .shared_arith = "off";

dffeas \mif_next_offset[27] (
	.clk(clk),
	.d(\Add1~109_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[27]~q ),
	.prn(vcc));
defparam \mif_next_offset[27] .is_wysiwyg = "true";
defparam \mif_next_offset[27] .power_up = "low";

cyclonev_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[27]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_27),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(\Add0~110 ),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

cyclonev_lcell_comb \Add1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~113_sumout ),
	.cout(\Add1~114 ),
	.shareout());
defparam \Add1~113 .extended_lut = "off";
defparam \Add1~113 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~113 .shared_arith = "off";

dffeas \mif_next_offset[28] (
	.clk(clk),
	.d(\Add1~113_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[28]~q ),
	.prn(vcc));
defparam \mif_next_offset[28] .is_wysiwyg = "true";
defparam \mif_next_offset[28] .power_up = "low";

cyclonev_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[28]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_28),
	.datag(gnd),
	.cin(\Add0~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

cyclonev_lcell_comb \Add1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~117_sumout ),
	.cout(\Add1~118 ),
	.shareout());
defparam \Add1~117 .extended_lut = "off";
defparam \Add1~117 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~117 .shared_arith = "off";

dffeas \mif_next_offset[29] (
	.clk(clk),
	.d(\Add1~117_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[29]~q ),
	.prn(vcc));
defparam \mif_next_offset[29] .is_wysiwyg = "true";
defparam \mif_next_offset[29] .power_up = "low";

cyclonev_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[29]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_29),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

cyclonev_lcell_comb \Add1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~121_sumout ),
	.cout(\Add1~122 ),
	.shareout());
defparam \Add1~121 .extended_lut = "off";
defparam \Add1~121 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~121 .shared_arith = "off";

dffeas \mif_next_offset[30] (
	.clk(clk),
	.d(\Add1~121_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[30]~q ),
	.prn(vcc));
defparam \mif_next_offset[30] .is_wysiwyg = "true";
defparam \mif_next_offset[30] .power_up = "low";

cyclonev_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[30]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_30),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

cyclonev_lcell_comb \Add1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~125_sumout ),
	.cout(),
	.shareout());
defparam \Add1~125 .extended_lut = "off";
defparam \Add1~125 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~125 .shared_arith = "off";

dffeas \mif_next_offset[31] (
	.clk(clk),
	.d(\Add1~125_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mif_next_offset~0_combout ),
	.sload(gnd),
	.ena(\mif_next_offset[28]~1_combout ),
	.q(\mif_next_offset[31]~q ),
	.prn(vcc));
defparam \mif_next_offset[31] .is_wysiwyg = "true";
defparam \mif_next_offset[31] .power_up = "low";

cyclonev_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\mif_next_offset[31]~q ),
	.datae(gnd),
	.dataf(!mif_base_addr_31),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h00000000000000FF;
defparam \Add3~17 .shared_arith = "off";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~13 .shared_arith = "off";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~9 .shared_arith = "off";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~21 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \av_mif_addr[2]~0 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\mif_len_cnt[1]~q ),
	.datac(!\mif_rec_len[1]~q ),
	.datad(!\mif_rec_len[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_mif_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_mif_addr[2]~0 .extended_lut = "off";
defparam \av_mif_addr[2]~0 .lut_mask = 64'h8241824182418241;
defparam \av_mif_addr[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \av_mif_addr[2]~1 (
	.dataa(!\mif_len_cnt[4]~q ),
	.datab(!\mif_len_cnt[3]~q ),
	.datac(!\mif_rec_len[4]~q ),
	.datad(!\mif_rec_len[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_mif_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_mif_addr[2]~1 .extended_lut = "off";
defparam \av_mif_addr[2]~1 .lut_mask = 64'h8421842184218421;
defparam \av_mif_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \av_mif_addr[2]~2 (
	.dataa(!\mif_len_cnt[2]~q ),
	.datab(!\mif_rec_len[2]~q ),
	.datac(!\av_mif_addr[2]~0_combout ),
	.datad(!\av_mif_addr[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_mif_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_mif_addr[2]~2 .extended_lut = "off";
defparam \av_mif_addr[2]~2 .lut_mask = 64'h0009000900090009;
defparam \av_mif_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \av_mif_addr[2]~3 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!\Selector2~1_combout ),
	.datad(!\mif_rec_data~0_combout ),
	.datae(!\av_mif_addr[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_mif_addr[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_mif_addr[2]~3 .extended_lut = "off";
defparam \av_mif_addr[2]~3 .lut_mask = 64'h0F7F0F0F0F7F0F0F;
defparam \av_mif_addr[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout());
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~41 .shared_arith = "off";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout());
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~37 .shared_arith = "off";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~25 .shared_arith = "off";

dffeas \mif_rec_addr[8] (
	.clk(clk),
	.d(stream_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[8]~q ),
	.prn(vcc));
defparam \mif_rec_addr[8] .is_wysiwyg = "true";
defparam \mif_rec_addr[8] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~29 .shared_arith = "off";

dffeas \mif_rec_addr[9] (
	.clk(clk),
	.d(stream_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[9]~q ),
	.prn(vcc));
defparam \mif_rec_addr[9] .is_wysiwyg = "true";
defparam \mif_rec_addr[9] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!av_mif_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~33 .shared_arith = "off";

dffeas \mif_rec_addr[10] (
	.clk(clk),
	.d(stream_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_next_state.AV_DEC_HDR~0_combout ),
	.q(\mif_rec_addr[10]~q ),
	.prn(vcc));
defparam \mif_rec_addr[10] .is_wysiwyg = "true";
defparam \mif_rec_addr[10] .power_up = "low";

cyclonev_lcell_comb \stream_read~0 (
	.dataa(!\Selector1~2_combout ),
	.datab(!\Selector2~3_combout ),
	.datac(!\Selector1~4_combout ),
	.datad(!\Selector1~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stream_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stream_read~0 .extended_lut = "off";
defparam \stream_read~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \stream_read~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ctrl_req~0 (
	.dataa(!\mif_len_cnt[0]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!av_ctrl_req1),
	.datad(!ctrl_op_done),
	.datae(!\mif_rec_data~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ctrl_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ctrl_req~0 .extended_lut = "off";
defparam \av_ctrl_req~0 .lut_mask = 64'h0F007F770F007F77;
defparam \av_ctrl_req~0 .shared_arith = "off";

cyclonev_lcell_comb \pll_go~0 (
	.dataa(!\av_state.AV_DEC_HDR~q ),
	.datab(!\Equal2~0_combout ),
	.datac(!\invalid_rec~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_go~0 .extended_lut = "off";
defparam \pll_go~0 .lut_mask = 64'h0101010101010101;
defparam \pll_go~0 .shared_arith = "off";

cyclonev_lcell_comb \always6~0 (
	.dataa(!stream_address_14),
	.datab(!stream_address_15),
	.datac(!stream_address_16),
	.datad(!mif_base_addr_14),
	.datae(!mif_base_addr_15),
	.dataf(!mif_base_addr_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'h8040201008040201;
defparam \always6~0 .shared_arith = "off";

cyclonev_lcell_comb \always6~1 (
	.dataa(!stream_address_26),
	.datab(!stream_address_27),
	.datac(!stream_address_28),
	.datad(!mif_base_addr_26),
	.datae(!mif_base_addr_27),
	.dataf(!mif_base_addr_28),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~1 .extended_lut = "off";
defparam \always6~1 .lut_mask = 64'h8040201008040201;
defparam \always6~1 .shared_arith = "off";

cyclonev_lcell_comb \always6~2 (
	.dataa(!stream_address_29),
	.datab(!stream_address_30),
	.datac(!stream_address_31),
	.datad(!mif_base_addr_29),
	.datae(!mif_base_addr_30),
	.dataf(!mif_base_addr_31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~2 .extended_lut = "off";
defparam \always6~2 .lut_mask = 64'h8040201008040201;
defparam \always6~2 .shared_arith = "off";

cyclonev_lcell_comb \always6~3 (
	.dataa(!stream_address_0),
	.datab(!stream_address_1),
	.datac(!stream_read1),
	.datad(!mif_base_addr_0),
	.datae(!reconfig_mif_waitrequest),
	.dataf(!mif_base_addr_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~3 .extended_lut = "off";
defparam \always6~3 .lut_mask = 64'h0804000002010000;
defparam \always6~3 .shared_arith = "off";

cyclonev_lcell_comb \always6~4 (
	.dataa(!stream_address_2),
	.datab(!stream_address_3),
	.datac(!stream_address_4),
	.datad(!mif_base_addr_2),
	.datae(!mif_base_addr_3),
	.dataf(!mif_base_addr_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~4 .extended_lut = "off";
defparam \always6~4 .lut_mask = 64'h8040201008040201;
defparam \always6~4 .shared_arith = "off";

cyclonev_lcell_comb \always6~5 (
	.dataa(!stream_address_5),
	.datab(!stream_address_6),
	.datac(!stream_address_7),
	.datad(!mif_base_addr_5),
	.datae(!mif_base_addr_6),
	.dataf(!mif_base_addr_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~5 .extended_lut = "off";
defparam \always6~5 .lut_mask = 64'h8040201008040201;
defparam \always6~5 .shared_arith = "off";

cyclonev_lcell_comb \always6~6 (
	.dataa(!stream_address_8),
	.datab(!stream_address_9),
	.datac(!stream_address_10),
	.datad(!mif_base_addr_8),
	.datae(!mif_base_addr_9),
	.dataf(!mif_base_addr_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~6 .extended_lut = "off";
defparam \always6~6 .lut_mask = 64'h8040201008040201;
defparam \always6~6 .shared_arith = "off";

cyclonev_lcell_comb \always6~7 (
	.dataa(!stream_address_11),
	.datab(!stream_address_12),
	.datac(!stream_address_13),
	.datad(!mif_base_addr_11),
	.datae(!mif_base_addr_12),
	.dataf(!mif_base_addr_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~7 .extended_lut = "off";
defparam \always6~7 .lut_mask = 64'h8040201008040201;
defparam \always6~7 .shared_arith = "off";

cyclonev_lcell_comb \always6~8 (
	.dataa(!\always6~3_combout ),
	.datab(!\always6~4_combout ),
	.datac(!\always6~5_combout ),
	.datad(!\always6~6_combout ),
	.datae(!\always6~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~8 .extended_lut = "off";
defparam \always6~8 .lut_mask = 64'h0000000100000001;
defparam \always6~8 .shared_arith = "off";

cyclonev_lcell_comb \always6~9 (
	.dataa(!stream_address_17),
	.datab(!stream_address_18),
	.datac(!stream_address_19),
	.datad(!mif_base_addr_17),
	.datae(!mif_base_addr_18),
	.dataf(!mif_base_addr_19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~9 .extended_lut = "off";
defparam \always6~9 .lut_mask = 64'h8040201008040201;
defparam \always6~9 .shared_arith = "off";

cyclonev_lcell_comb \always6~10 (
	.dataa(!stream_address_20),
	.datab(!stream_address_21),
	.datac(!mif_base_addr_20),
	.datad(!mif_base_addr_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~10 .extended_lut = "off";
defparam \always6~10 .lut_mask = 64'h8421842184218421;
defparam \always6~10 .shared_arith = "off";

cyclonev_lcell_comb \always6~11 (
	.dataa(!stream_address_23),
	.datab(!stream_address_24),
	.datac(!stream_address_25),
	.datad(!mif_base_addr_23),
	.datae(!mif_base_addr_24),
	.dataf(!mif_base_addr_25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~11 .extended_lut = "off";
defparam \always6~11 .lut_mask = 64'h8040201008040201;
defparam \always6~11 .shared_arith = "off";

cyclonev_lcell_comb \always6~12 (
	.dataa(!stream_address_22),
	.datab(!mif_base_addr_22),
	.datac(!\always6~9_combout ),
	.datad(!\always6~10_combout ),
	.datae(!\always6~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~12 .extended_lut = "off";
defparam \always6~12 .lut_mask = 64'h0000000900000009;
defparam \always6~12 .shared_arith = "off";

cyclonev_lcell_comb \always6~13 (
	.dataa(!\always6~0_combout ),
	.datab(!\always6~1_combout ),
	.datac(!\always6~2_combout ),
	.datad(!\always6~8_combout ),
	.datae(!\always6~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~13 .extended_lut = "off";
defparam \always6~13 .lut_mask = 64'h0000000100000001;
defparam \always6~13 .shared_arith = "off";

dffeas first_mif_entry(
	.clk(clk),
	.d(\always6~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\first_mif_entry~q ),
	.prn(vcc));
defparam first_mif_entry.is_wysiwyg = "true";
defparam first_mif_entry.power_up = "low";

cyclonev_lcell_comb \av_opcode_err~0 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\av_state.AV_IDLE~q ),
	.datac(!\rec_is_som~0_combout ),
	.datad(!\mif_strm_active~q ),
	.datae(!\invalid_rec~1_combout ),
	.dataf(!\first_mif_entry~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_opcode_err~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_opcode_err~0 .extended_lut = "off";
defparam \av_opcode_err~0 .lut_mask = 64'h00550044F0F5F0F4;
defparam \av_opcode_err~0 .shared_arith = "off";

cyclonev_lcell_comb \av_done~0 (
	.dataa(!\av_state.AV_IDLE~q ),
	.datab(!\Selector0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_done~0 .extended_lut = "off";
defparam \av_done~0 .lut_mask = 64'h4444444444444444;
defparam \av_done~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!\mif_rec_addr[2]~q ),
	.datab(!\mif_rec_addr[1]~q ),
	.datac(!\mif_rec_addr[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'h4040404040404040;
defparam \Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb rec_is_cgb(
	.dataa(!\Equal2~0_combout ),
	.datab(!\av_state.AV_IDLE~q ),
	.datac(!\mif_rec_addr[4]~q ),
	.datad(!\mif_rec_addr[3]~q ),
	.datae(!\Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rec_is_cgb~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam rec_is_cgb.extended_lut = "off";
defparam rec_is_cgb.lut_mask = 64'h0000100000001000;
defparam rec_is_cgb.shared_arith = "off";

cyclonev_lcell_comb \rec_is_type~0 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\av_state.AV_IDLE~q ),
	.datac(!\mif_rec_addr[1]~q ),
	.datad(!\mif_rec_addr[0]~q ),
	.datae(!\Equal6~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rec_is_type~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rec_is_type~0 .extended_lut = "off";
defparam \rec_is_type~0 .lut_mask = 64'h0000010000000100;
defparam \rec_is_type~0 .shared_arith = "off";

cyclonev_lcell_comb \av_mif_type~0 (
	.dataa(!mif_rec_addr_6),
	.datab(!\rec_is_type~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_mif_type~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_mif_type~0 .extended_lut = "off";
defparam \av_mif_type~0 .lut_mask = 64'h1111111111111111;
defparam \av_mif_type~0 .shared_arith = "off";

cyclonev_lcell_comb \av_mif_type~1 (
	.dataa(!mif_rec_addr_5),
	.datab(!\rec_is_type~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_mif_type~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_mif_type~1 .extended_lut = "off";
defparam \av_mif_type~1 .lut_mask = 64'h1111111111111111;
defparam \av_mif_type~1 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_av_xcvr_reconfig_mif_ctrl (
	uif_rdata_5,
	uif_rdata_6,
	uif_rdata_7,
	uif_rdata_8,
	uif_rdata_9,
	uif_rdata_10,
	uif_rdata_11,
	uif_rdata_12,
	uif_rdata_13,
	uif_rdata_14,
	uif_rdata_15,
	uif_rdata_16,
	uif_rdata_17,
	uif_rdata_18,
	uif_rdata_19,
	uif_rdata_20,
	uif_rdata_21,
	uif_rdata_22,
	uif_rdata_23,
	uif_rdata_24,
	uif_rdata_25,
	uif_rdata_26,
	uif_rdata_27,
	uif_rdata_28,
	uif_rdata_29,
	uif_rdata_30,
	uif_rdata_31,
	ctrl_addr_1,
	ctrl_addr_2,
	ctrl_addr_0,
	av_mif_addr_4,
	av_mif_addr_5,
	av_mif_addr_2,
	av_mif_addr_1,
	av_mif_addr_0,
	av_mif_addr_3,
	av_mif_addr_8,
	av_mif_addr_9,
	av_mif_addr_10,
	av_mif_addr_7,
	av_mif_addr_6,
	ctrl_addr_4,
	ctrl_addr_5,
	ctrl_addr_6,
	ctrl_addr_7,
	ctrl_addr_8,
	ctrl_addr_9,
	ctrl_addr_10,
	uif_busy1,
	reset,
	uif_writedata_0,
	uif_mode_1,
	uif_mode_0,
	Equal5,
	uif_rdata_0,
	uif_addr_offset_0,
	uif_writedata_1,
	uif_rdata_1,
	uif_addr_offset_1,
	uif_writedata_2,
	uif_ctrl_0,
	uif_addr_offset_2,
	uif_rdata_2,
	uif_writedata_3,
	uif_ctrl_1,
	uif_addr_offset_3,
	uif_rdata_3,
	uif_writedata_4,
	uif_rdata_4,
	uif_addr_offset_4,
	uif_writedata_5,
	uif_addr_offset_5,
	uif_writedata_6,
	uif_addr_offset_6,
	uif_writedata_7,
	uif_addr_offset_7,
	uif_writedata_8,
	uif_addr_offset_8,
	uif_writedata_9,
	uif_addr_err1,
	uif_addr_offset_9,
	uif_writedata_10,
	uif_addr_offset_10,
	uif_writedata_11,
	uif_addr_offset_11,
	uif_writedata_12,
	uif_writedata_13,
	uif_writedata_14,
	uif_writedata_15,
	uif_writedata_16,
	uif_writedata_17,
	uif_writedata_18,
	uif_writedata_19,
	uif_writedata_20,
	uif_writedata_21,
	uif_writedata_22,
	uif_writedata_23,
	uif_writedata_24,
	uif_writedata_25,
	uif_writedata_26,
	uif_writedata_27,
	uif_writedata_28,
	uif_writedata_29,
	uif_writedata_30,
	uif_writedata_31,
	ctrl_opcode_1,
	ctrl_opcode_2,
	ctrl_opcode_0,
	ctrl_go1,
	ctrl_lock1,
	av_ctrl_req,
	waitrequest_to_ctrl,
	ctrl_op_done,
	mif_err_reg_4,
	mif_err_reg_1,
	mif_err_reg_0,
	ctrl_av_go1,
	ctrl_rdata,
	uif_go,
	mif_base_addr_0,
	mif_base_addr_1,
	mif_base_addr_2,
	mif_base_addr_3,
	mif_base_addr_4,
	mif_base_addr_5,
	mif_base_addr_6,
	mif_base_addr_7,
	mif_base_addr_8,
	mif_base_addr_9,
	mif_base_addr_10,
	mif_base_addr_11,
	mif_base_addr_12,
	mif_base_addr_13,
	mif_base_addr_14,
	mif_base_addr_15,
	mif_base_addr_16,
	readdata_for_user_16,
	mif_base_addr_17,
	readdata_for_user_17,
	mif_base_addr_18,
	readdata_for_user_18,
	mif_base_addr_19,
	readdata_for_user_19,
	mif_base_addr_20,
	readdata_for_user_20,
	mif_base_addr_21,
	readdata_for_user_21,
	mif_base_addr_22,
	readdata_for_user_22,
	mif_base_addr_23,
	readdata_for_user_23,
	mif_base_addr_24,
	readdata_for_user_24,
	mif_base_addr_25,
	readdata_for_user_25,
	mif_base_addr_26,
	readdata_for_user_26,
	mif_base_addr_27,
	readdata_for_user_27,
	mif_base_addr_28,
	readdata_for_user_28,
	mif_base_addr_29,
	readdata_for_user_29,
	mif_base_addr_30,
	readdata_for_user_30,
	mif_base_addr_31,
	readdata_for_user_31,
	av_addr_burst,
	ctrl_wdata_1,
	ctrl_wdata_2,
	ctrl_wdata_0,
	ctrl_wdata_3,
	ctrl_addr_3,
	av_opcode_err,
	ctrl_wdata_4,
	ctrl_wdata_5,
	ctrl_wdata_6,
	ctrl_wdata_7,
	ctrl_wdata_8,
	ctrl_wdata_9,
	ctrl_wdata_10,
	ctrl_wdata_11,
	ctrl_addr_11,
	ctrl_wdata_12,
	ctrl_wdata_13,
	ctrl_wdata_14,
	ctrl_wdata_15,
	av_done,
	mif_rec_data_1,
	mif_rec_data_2,
	mif_rec_data_0,
	mif_rec_data_3,
	av_mif_type_valid,
	av_mif_type_1,
	av_mif_type_0,
	mif_rec_data_4,
	mif_rec_data_5,
	mif_rec_data_6,
	mif_rec_data_7,
	mif_rec_data_8,
	mif_rec_data_9,
	mif_rec_data_10,
	mif_rec_data_11,
	mif_rec_data_12,
	mif_rec_data_13,
	mif_rec_data_14,
	mif_rec_data_15,
	mif_addr_mode1,
	clk)/* synthesis synthesis_greybox=0 */;
output 	uif_rdata_5;
output 	uif_rdata_6;
output 	uif_rdata_7;
output 	uif_rdata_8;
output 	uif_rdata_9;
output 	uif_rdata_10;
output 	uif_rdata_11;
output 	uif_rdata_12;
output 	uif_rdata_13;
output 	uif_rdata_14;
output 	uif_rdata_15;
output 	uif_rdata_16;
output 	uif_rdata_17;
output 	uif_rdata_18;
output 	uif_rdata_19;
output 	uif_rdata_20;
output 	uif_rdata_21;
output 	uif_rdata_22;
output 	uif_rdata_23;
output 	uif_rdata_24;
output 	uif_rdata_25;
output 	uif_rdata_26;
output 	uif_rdata_27;
output 	uif_rdata_28;
output 	uif_rdata_29;
output 	uif_rdata_30;
output 	uif_rdata_31;
output 	ctrl_addr_1;
output 	ctrl_addr_2;
output 	ctrl_addr_0;
input 	av_mif_addr_4;
input 	av_mif_addr_5;
input 	av_mif_addr_2;
input 	av_mif_addr_1;
input 	av_mif_addr_0;
input 	av_mif_addr_3;
input 	av_mif_addr_8;
input 	av_mif_addr_9;
input 	av_mif_addr_10;
input 	av_mif_addr_7;
input 	av_mif_addr_6;
output 	ctrl_addr_4;
output 	ctrl_addr_5;
output 	ctrl_addr_6;
output 	ctrl_addr_7;
output 	ctrl_addr_8;
output 	ctrl_addr_9;
output 	ctrl_addr_10;
output 	uif_busy1;
input 	reset;
input 	uif_writedata_0;
input 	uif_mode_1;
input 	uif_mode_0;
output 	Equal5;
output 	uif_rdata_0;
input 	uif_addr_offset_0;
input 	uif_writedata_1;
output 	uif_rdata_1;
input 	uif_addr_offset_1;
input 	uif_writedata_2;
input 	uif_ctrl_0;
input 	uif_addr_offset_2;
output 	uif_rdata_2;
input 	uif_writedata_3;
input 	uif_ctrl_1;
input 	uif_addr_offset_3;
output 	uif_rdata_3;
input 	uif_writedata_4;
output 	uif_rdata_4;
input 	uif_addr_offset_4;
input 	uif_writedata_5;
input 	uif_addr_offset_5;
input 	uif_writedata_6;
input 	uif_addr_offset_6;
input 	uif_writedata_7;
input 	uif_addr_offset_7;
input 	uif_writedata_8;
input 	uif_addr_offset_8;
input 	uif_writedata_9;
output 	uif_addr_err1;
input 	uif_addr_offset_9;
input 	uif_writedata_10;
input 	uif_addr_offset_10;
input 	uif_writedata_11;
input 	uif_addr_offset_11;
input 	uif_writedata_12;
input 	uif_writedata_13;
input 	uif_writedata_14;
input 	uif_writedata_15;
input 	uif_writedata_16;
input 	uif_writedata_17;
input 	uif_writedata_18;
input 	uif_writedata_19;
input 	uif_writedata_20;
input 	uif_writedata_21;
input 	uif_writedata_22;
input 	uif_writedata_23;
input 	uif_writedata_24;
input 	uif_writedata_25;
input 	uif_writedata_26;
input 	uif_writedata_27;
input 	uif_writedata_28;
input 	uif_writedata_29;
input 	uif_writedata_30;
input 	uif_writedata_31;
output 	ctrl_opcode_1;
output 	ctrl_opcode_2;
output 	ctrl_opcode_0;
output 	ctrl_go1;
output 	ctrl_lock1;
input 	av_ctrl_req;
input 	waitrequest_to_ctrl;
output 	ctrl_op_done;
output 	mif_err_reg_4;
output 	mif_err_reg_1;
output 	mif_err_reg_0;
output 	ctrl_av_go1;
input 	[31:0] ctrl_rdata;
input 	uif_go;
output 	mif_base_addr_0;
output 	mif_base_addr_1;
output 	mif_base_addr_2;
output 	mif_base_addr_3;
output 	mif_base_addr_4;
output 	mif_base_addr_5;
output 	mif_base_addr_6;
output 	mif_base_addr_7;
output 	mif_base_addr_8;
output 	mif_base_addr_9;
output 	mif_base_addr_10;
output 	mif_base_addr_11;
output 	mif_base_addr_12;
output 	mif_base_addr_13;
output 	mif_base_addr_14;
output 	mif_base_addr_15;
output 	mif_base_addr_16;
input 	readdata_for_user_16;
output 	mif_base_addr_17;
input 	readdata_for_user_17;
output 	mif_base_addr_18;
input 	readdata_for_user_18;
output 	mif_base_addr_19;
input 	readdata_for_user_19;
output 	mif_base_addr_20;
input 	readdata_for_user_20;
output 	mif_base_addr_21;
input 	readdata_for_user_21;
output 	mif_base_addr_22;
input 	readdata_for_user_22;
output 	mif_base_addr_23;
input 	readdata_for_user_23;
output 	mif_base_addr_24;
input 	readdata_for_user_24;
output 	mif_base_addr_25;
input 	readdata_for_user_25;
output 	mif_base_addr_26;
input 	readdata_for_user_26;
output 	mif_base_addr_27;
input 	readdata_for_user_27;
output 	mif_base_addr_28;
input 	readdata_for_user_28;
output 	mif_base_addr_29;
input 	readdata_for_user_29;
output 	mif_base_addr_30;
input 	readdata_for_user_30;
output 	mif_base_addr_31;
input 	readdata_for_user_31;
input 	av_addr_burst;
output 	ctrl_wdata_1;
output 	ctrl_wdata_2;
output 	ctrl_wdata_0;
output 	ctrl_wdata_3;
output 	ctrl_addr_3;
input 	av_opcode_err;
output 	ctrl_wdata_4;
output 	ctrl_wdata_5;
output 	ctrl_wdata_6;
output 	ctrl_wdata_7;
output 	ctrl_wdata_8;
output 	ctrl_wdata_9;
output 	ctrl_wdata_10;
output 	ctrl_wdata_11;
output 	ctrl_addr_11;
output 	ctrl_wdata_12;
output 	ctrl_wdata_13;
output 	ctrl_wdata_14;
output 	ctrl_wdata_15;
input 	av_done;
input 	mif_rec_data_1;
input 	mif_rec_data_2;
input 	mif_rec_data_0;
input 	mif_rec_data_3;
input 	av_mif_type_valid;
input 	av_mif_type_1;
input 	av_mif_type_0;
input 	mif_rec_data_4;
input 	mif_rec_data_5;
input 	mif_rec_data_6;
input 	mif_rec_data_7;
input 	mif_rec_data_8;
input 	mif_rec_data_9;
input 	mif_rec_data_10;
input 	mif_rec_data_11;
input 	mif_rec_data_12;
input 	mif_rec_data_13;
input 	mif_rec_data_14;
input 	mif_rec_data_15;
output 	mif_addr_mode1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ctrl_wdata~0_combout ;
wire \always1~0_combout ;
wire \Equal3~0_combout ;
wire \uif_rdata[11]~3_combout ;
wire \uif_rdata[2]~0_combout ;
wire \always0~0_combout ;
wire \mif_strm_start~0_combout ;
wire \mif_strm_start~1_combout ;
wire \mif_strm_start~q ;
wire \ctrl_next_state~0_combout ;
wire \set_uif_ctrl_req~0_combout ;
wire \uif_ctrl_req~0_combout ;
wire \uif_ctrl_req~q ;
wire \chn_chk_active~0_combout ;
wire \chn_chk_active~q ;
wire \always3~0_combout ;
wire \Selector8~0_combout ;
wire \ctrl_state.CTRL_WF_AV~q ;
wire \Selector10~0_combout ;
wire \Selector10~1_combout ;
wire \ctrl_state.CTRL_CHK_ADDR~q ;
wire \Selector6~0_combout ;
wire \ctrl_state.CTRL_MIF_WR~q ;
wire \Selector9~0_combout ;
wire \ctrl_state.CTRL_MIF_RD~q ;
wire \ctrl_state.CTRL_CHK_CHN~q ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \ctrl_state.CTRL_WF_B~q ;
wire \Selector5~1_combout ;
wire \ctrl_next_state.CTRL_RMW~0_combout ;
wire \ctrl_state.CTRL_RMW~q ;
wire \av_ctrl_req_dly~q ;
wire \always9~0_combout ;
wire \mux_mif_addr[4]~0_combout ;
wire \mux_mif_addr[5]~1_combout ;
wire \mux_mif_addr[2]~2_combout ;
wire \mux_mif_addr[1]~3_combout ;
wire \mux_mif_addr[0]~4_combout ;
wire \mux_mif_addr[3]~5_combout ;
wire \Equal14~0_combout ;
wire \Equal14~1_combout ;
wire \Equal14~2_combout ;
wire \Equal14~3_combout ;
wire \Equal22~0_combout ;
wire \Equal22~1_combout ;
wire \Equal17~0_combout ;
wire \Equal17~1_combout ;
wire \ctrl_wdata~1_combout ;
wire \Equal14~4_combout ;
wire \Equal14~5_combout ;
wire \Equal15~0_combout ;
wire \mux_mif_addr[6]~6_combout ;
wire \Equal23~0_combout ;
wire \Equal23~1_combout ;
wire \WideNor1~0_combout ;
wire \rmw_offset~0_combout ;
wire \rmw_offset~q ;
wire \ctrl_next_state~1_combout ;
wire \Selector5~2_combout ;
wire \Selector5~3_combout ;
wire \ctrl_state.CTRL_IDLE~q ;
wire \ctrl_next_state.CTRL_CHK_CHN~0_combout ;
wire \always6~0_combout ;
wire \ctrl_addr[1]~0_combout ;
wire \uif_rdata~12_combout ;
wire \uif_rdata~8_combout ;
wire \uif_rdata~1_combout ;
wire \uif_rdata~2_combout ;
wire \uif_rdata~4_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \uif_addr_err_d~combout ;
wire \ctrl_opcode~0_combout ;
wire \ctrl_opcode~1_combout ;
wire \ctrl_opcode[1]~2_combout ;
wire \ctrl_opcode~3_combout ;
wire \ctrl_opcode~4_combout ;
wire \ctrl_lock~0_combout ;
wire \mif_clr_error~0_combout ;
wire \mif_clr_error~q ;
wire \channel_id~2_combout ;
wire \always7~0_combout ;
wire \channel_id[0]~1_combout ;
wire \channel_id[0]~q ;
wire \channel_id~0_combout ;
wire \channel_id[1]~q ;
wire \channel_id~3_combout ;
wire \channel_id[3]~q ;
wire \channel_id~4_combout ;
wire \channel_id[2]~q ;
wire \av_chn_mismatch~0_combout ;
wire \av_chn_mismatch~1_combout ;
wire \av_chn_mismatch~q ;
wire \mif_err_reg~0_combout ;
wire \mif_err_reg~1_combout ;
wire \mif_err_reg~2_combout ;
wire \ctrl_av_go~0_combout ;
wire \mif_base_addr[31]~0_combout ;
wire \WideOr16~0_combout ;
wire \saved_read_data[1]~q ;
wire \ctrl_wdata~2_combout ;
wire \Equal23~2_combout ;
wire \saved_read_data[2]~q ;
wire \ctrl_wdata~3_combout ;
wire \ctrl_wdata~4_combout ;
wire \saved_read_data[0]~q ;
wire \ctrl_wdata~5_combout ;
wire \saved_read_data[3]~q ;
wire \WideOr14~0_combout ;
wire \ctrl_wdata~6_combout ;
wire \ctrl_addr~1_combout ;
wire \ctrl_addr~2_combout ;
wire \saved_read_data[4]~q ;
wire \ctrl_wdata~7_combout ;
wire \WideOr14~combout ;
wire \saved_read_data[5]~q ;
wire \ctrl_wdata~8_combout ;
wire \saved_read_data[6]~q ;
wire \Equal20~0_combout ;
wire \ctrl_wdata[6]~9_combout ;
wire \ctrl_wdata~10_combout ;
wire \saved_read_data[7]~q ;
wire \ctrl_wdata~11_combout ;
wire \ctrl_wdata~12_combout ;
wire \saved_read_data[8]~q ;
wire \ctrl_wdata~13_combout ;
wire \ctrl_wdata~14_combout ;
wire \saved_read_data[9]~q ;
wire \ctrl_wdata~15_combout ;
wire \ctrl_wdata~16_combout ;
wire \saved_read_data[10]~q ;
wire \ctrl_wdata~17_combout ;
wire \ctrl_wdata~18_combout ;
wire \saved_read_data[11]~q ;
wire \ctrl_wdata~19_combout ;
wire \ctrl_wdata~20_combout ;
wire \ctrl_addr~3_combout ;
wire \saved_read_data[12]~q ;
wire \ctrl_wdata~21_combout ;
wire \ctrl_wdata~22_combout ;
wire \Equal16~0_combout ;
wire \saved_read_data[13]~q ;
wire \ctrl_wdata~23_combout ;
wire \ctrl_wdata~24_combout ;
wire \saved_read_data[14]~q ;
wire \ctrl_wdata~25_combout ;
wire \ctrl_wdata~26_combout ;
wire \saved_read_data[15]~q ;
wire \ctrl_wdata~27_combout ;
wire \ctrl_wdata~28_combout ;
wire \mif_addr_mode~0_combout ;


dffeas \uif_rdata[5] (
	.clk(clk),
	.d(mif_base_addr_5),
	.asdata(ctrl_rdata[5]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_5),
	.prn(vcc));
defparam \uif_rdata[5] .is_wysiwyg = "true";
defparam \uif_rdata[5] .power_up = "low";

dffeas \uif_rdata[6] (
	.clk(clk),
	.d(mif_base_addr_6),
	.asdata(ctrl_rdata[6]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_6),
	.prn(vcc));
defparam \uif_rdata[6] .is_wysiwyg = "true";
defparam \uif_rdata[6] .power_up = "low";

dffeas \uif_rdata[7] (
	.clk(clk),
	.d(mif_base_addr_7),
	.asdata(ctrl_rdata[7]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_7),
	.prn(vcc));
defparam \uif_rdata[7] .is_wysiwyg = "true";
defparam \uif_rdata[7] .power_up = "low";

dffeas \uif_rdata[8] (
	.clk(clk),
	.d(mif_base_addr_8),
	.asdata(ctrl_rdata[8]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_8),
	.prn(vcc));
defparam \uif_rdata[8] .is_wysiwyg = "true";
defparam \uif_rdata[8] .power_up = "low";

dffeas \uif_rdata[9] (
	.clk(clk),
	.d(mif_base_addr_9),
	.asdata(ctrl_rdata[9]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_9),
	.prn(vcc));
defparam \uif_rdata[9] .is_wysiwyg = "true";
defparam \uif_rdata[9] .power_up = "low";

dffeas \uif_rdata[10] (
	.clk(clk),
	.d(mif_base_addr_10),
	.asdata(ctrl_rdata[10]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_10),
	.prn(vcc));
defparam \uif_rdata[10] .is_wysiwyg = "true";
defparam \uif_rdata[10] .power_up = "low";

dffeas \uif_rdata[11] (
	.clk(clk),
	.d(mif_base_addr_11),
	.asdata(ctrl_rdata[11]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_11),
	.prn(vcc));
defparam \uif_rdata[11] .is_wysiwyg = "true";
defparam \uif_rdata[11] .power_up = "low";

dffeas \uif_rdata[12] (
	.clk(clk),
	.d(mif_base_addr_12),
	.asdata(ctrl_rdata[12]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_12),
	.prn(vcc));
defparam \uif_rdata[12] .is_wysiwyg = "true";
defparam \uif_rdata[12] .power_up = "low";

dffeas \uif_rdata[13] (
	.clk(clk),
	.d(mif_base_addr_13),
	.asdata(ctrl_rdata[13]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_13),
	.prn(vcc));
defparam \uif_rdata[13] .is_wysiwyg = "true";
defparam \uif_rdata[13] .power_up = "low";

dffeas \uif_rdata[14] (
	.clk(clk),
	.d(mif_base_addr_14),
	.asdata(ctrl_rdata[14]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_14),
	.prn(vcc));
defparam \uif_rdata[14] .is_wysiwyg = "true";
defparam \uif_rdata[14] .power_up = "low";

dffeas \uif_rdata[15] (
	.clk(clk),
	.d(mif_base_addr_15),
	.asdata(ctrl_rdata[15]),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_15),
	.prn(vcc));
defparam \uif_rdata[15] .is_wysiwyg = "true";
defparam \uif_rdata[15] .power_up = "low";

dffeas \uif_rdata[16] (
	.clk(clk),
	.d(mif_base_addr_16),
	.asdata(readdata_for_user_16),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_16),
	.prn(vcc));
defparam \uif_rdata[16] .is_wysiwyg = "true";
defparam \uif_rdata[16] .power_up = "low";

dffeas \uif_rdata[17] (
	.clk(clk),
	.d(mif_base_addr_17),
	.asdata(readdata_for_user_17),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_17),
	.prn(vcc));
defparam \uif_rdata[17] .is_wysiwyg = "true";
defparam \uif_rdata[17] .power_up = "low";

dffeas \uif_rdata[18] (
	.clk(clk),
	.d(mif_base_addr_18),
	.asdata(readdata_for_user_18),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_18),
	.prn(vcc));
defparam \uif_rdata[18] .is_wysiwyg = "true";
defparam \uif_rdata[18] .power_up = "low";

dffeas \uif_rdata[19] (
	.clk(clk),
	.d(mif_base_addr_19),
	.asdata(readdata_for_user_19),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_19),
	.prn(vcc));
defparam \uif_rdata[19] .is_wysiwyg = "true";
defparam \uif_rdata[19] .power_up = "low";

dffeas \uif_rdata[20] (
	.clk(clk),
	.d(mif_base_addr_20),
	.asdata(readdata_for_user_20),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_20),
	.prn(vcc));
defparam \uif_rdata[20] .is_wysiwyg = "true";
defparam \uif_rdata[20] .power_up = "low";

dffeas \uif_rdata[21] (
	.clk(clk),
	.d(mif_base_addr_21),
	.asdata(readdata_for_user_21),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_21),
	.prn(vcc));
defparam \uif_rdata[21] .is_wysiwyg = "true";
defparam \uif_rdata[21] .power_up = "low";

dffeas \uif_rdata[22] (
	.clk(clk),
	.d(mif_base_addr_22),
	.asdata(readdata_for_user_22),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_22),
	.prn(vcc));
defparam \uif_rdata[22] .is_wysiwyg = "true";
defparam \uif_rdata[22] .power_up = "low";

dffeas \uif_rdata[23] (
	.clk(clk),
	.d(mif_base_addr_23),
	.asdata(readdata_for_user_23),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_23),
	.prn(vcc));
defparam \uif_rdata[23] .is_wysiwyg = "true";
defparam \uif_rdata[23] .power_up = "low";

dffeas \uif_rdata[24] (
	.clk(clk),
	.d(mif_base_addr_24),
	.asdata(readdata_for_user_24),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_24),
	.prn(vcc));
defparam \uif_rdata[24] .is_wysiwyg = "true";
defparam \uif_rdata[24] .power_up = "low";

dffeas \uif_rdata[25] (
	.clk(clk),
	.d(mif_base_addr_25),
	.asdata(readdata_for_user_25),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_25),
	.prn(vcc));
defparam \uif_rdata[25] .is_wysiwyg = "true";
defparam \uif_rdata[25] .power_up = "low";

dffeas \uif_rdata[26] (
	.clk(clk),
	.d(mif_base_addr_26),
	.asdata(readdata_for_user_26),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_26),
	.prn(vcc));
defparam \uif_rdata[26] .is_wysiwyg = "true";
defparam \uif_rdata[26] .power_up = "low";

dffeas \uif_rdata[27] (
	.clk(clk),
	.d(mif_base_addr_27),
	.asdata(readdata_for_user_27),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_27),
	.prn(vcc));
defparam \uif_rdata[27] .is_wysiwyg = "true";
defparam \uif_rdata[27] .power_up = "low";

dffeas \uif_rdata[28] (
	.clk(clk),
	.d(mif_base_addr_28),
	.asdata(readdata_for_user_28),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_28),
	.prn(vcc));
defparam \uif_rdata[28] .is_wysiwyg = "true";
defparam \uif_rdata[28] .power_up = "low";

dffeas \uif_rdata[29] (
	.clk(clk),
	.d(mif_base_addr_29),
	.asdata(readdata_for_user_29),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_29),
	.prn(vcc));
defparam \uif_rdata[29] .is_wysiwyg = "true";
defparam \uif_rdata[29] .power_up = "low";

dffeas \uif_rdata[30] (
	.clk(clk),
	.d(mif_base_addr_30),
	.asdata(readdata_for_user_30),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_30),
	.prn(vcc));
defparam \uif_rdata[30] .is_wysiwyg = "true";
defparam \uif_rdata[30] .power_up = "low";

dffeas \uif_rdata[31] (
	.clk(clk),
	.d(mif_base_addr_31),
	.asdata(readdata_for_user_31),
	.clrn(reset),
	.aload(gnd),
	.sclr(\uif_rdata[11]~3_combout ),
	.sload(!\always1~0_combout ),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_31),
	.prn(vcc));
defparam \uif_rdata[31] .is_wysiwyg = "true";
defparam \uif_rdata[31] .power_up = "low";

dffeas \ctrl_addr[1] (
	.clk(clk),
	.d(av_mif_addr_1),
	.asdata(uif_addr_offset_1),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_1),
	.prn(vcc));
defparam \ctrl_addr[1] .is_wysiwyg = "true";
defparam \ctrl_addr[1] .power_up = "low";

dffeas \ctrl_addr[2] (
	.clk(clk),
	.d(av_mif_addr_2),
	.asdata(uif_addr_offset_2),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_2),
	.prn(vcc));
defparam \ctrl_addr[2] .is_wysiwyg = "true";
defparam \ctrl_addr[2] .power_up = "low";

dffeas \ctrl_addr[0] (
	.clk(clk),
	.d(av_mif_addr_0),
	.asdata(uif_addr_offset_0),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_0),
	.prn(vcc));
defparam \ctrl_addr[0] .is_wysiwyg = "true";
defparam \ctrl_addr[0] .power_up = "low";

dffeas \ctrl_addr[4] (
	.clk(clk),
	.d(av_mif_addr_4),
	.asdata(uif_addr_offset_4),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_4),
	.prn(vcc));
defparam \ctrl_addr[4] .is_wysiwyg = "true";
defparam \ctrl_addr[4] .power_up = "low";

dffeas \ctrl_addr[5] (
	.clk(clk),
	.d(av_mif_addr_5),
	.asdata(uif_addr_offset_5),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_5),
	.prn(vcc));
defparam \ctrl_addr[5] .is_wysiwyg = "true";
defparam \ctrl_addr[5] .power_up = "low";

dffeas \ctrl_addr[6] (
	.clk(clk),
	.d(av_mif_addr_6),
	.asdata(uif_addr_offset_6),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_6),
	.prn(vcc));
defparam \ctrl_addr[6] .is_wysiwyg = "true";
defparam \ctrl_addr[6] .power_up = "low";

dffeas \ctrl_addr[7] (
	.clk(clk),
	.d(av_mif_addr_7),
	.asdata(uif_addr_offset_7),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_7),
	.prn(vcc));
defparam \ctrl_addr[7] .is_wysiwyg = "true";
defparam \ctrl_addr[7] .power_up = "low";

dffeas \ctrl_addr[8] (
	.clk(clk),
	.d(av_mif_addr_8),
	.asdata(uif_addr_offset_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_8),
	.prn(vcc));
defparam \ctrl_addr[8] .is_wysiwyg = "true";
defparam \ctrl_addr[8] .power_up = "low";

dffeas \ctrl_addr[9] (
	.clk(clk),
	.d(av_mif_addr_9),
	.asdata(uif_addr_offset_9),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_9),
	.prn(vcc));
defparam \ctrl_addr[9] .is_wysiwyg = "true";
defparam \ctrl_addr[9] .power_up = "low";

dffeas \ctrl_addr[10] (
	.clk(clk),
	.d(av_mif_addr_10),
	.asdata(uif_addr_offset_10),
	.clrn(reset),
	.aload(gnd),
	.sclr(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sload(\always6~0_combout ),
	.ena(\ctrl_addr[1]~0_combout ),
	.q(ctrl_addr_10),
	.prn(vcc));
defparam \ctrl_addr[10] .is_wysiwyg = "true";
defparam \ctrl_addr[10] .power_up = "low";

dffeas uif_busy(
	.clk(clk),
	.d(\ctrl_state.CTRL_IDLE~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_busy1),
	.prn(vcc));
defparam uif_busy.is_wysiwyg = "true";
defparam uif_busy.power_up = "low";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'h2222222222222222;
defparam \Equal5~0 .shared_arith = "off";

dffeas \uif_rdata[0] (
	.clk(clk),
	.d(\uif_rdata~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_0),
	.prn(vcc));
defparam \uif_rdata[0] .is_wysiwyg = "true";
defparam \uif_rdata[0] .power_up = "low";

dffeas \uif_rdata[1] (
	.clk(clk),
	.d(\uif_rdata~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_1),
	.prn(vcc));
defparam \uif_rdata[1] .is_wysiwyg = "true";
defparam \uif_rdata[1] .power_up = "low";

dffeas \uif_rdata[2] (
	.clk(clk),
	.d(\uif_rdata~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_2),
	.prn(vcc));
defparam \uif_rdata[2] .is_wysiwyg = "true";
defparam \uif_rdata[2] .power_up = "low";

dffeas \uif_rdata[3] (
	.clk(clk),
	.d(\uif_rdata~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_3),
	.prn(vcc));
defparam \uif_rdata[3] .is_wysiwyg = "true";
defparam \uif_rdata[3] .power_up = "low";

dffeas \uif_rdata[4] (
	.clk(clk),
	.d(\uif_rdata~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rdata[2]~0_combout ),
	.q(uif_rdata_4),
	.prn(vcc));
defparam \uif_rdata[4] .is_wysiwyg = "true";
defparam \uif_rdata[4] .power_up = "low";

dffeas uif_addr_err(
	.clk(clk),
	.d(\uif_addr_err_d~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_addr_err1),
	.prn(vcc));
defparam uif_addr_err.is_wysiwyg = "true";
defparam uif_addr_err.power_up = "low";

dffeas \ctrl_opcode[1] (
	.clk(clk),
	.d(\ctrl_opcode~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_opcode[1]~2_combout ),
	.q(ctrl_opcode_1),
	.prn(vcc));
defparam \ctrl_opcode[1] .is_wysiwyg = "true";
defparam \ctrl_opcode[1] .power_up = "low";

dffeas \ctrl_opcode[2] (
	.clk(clk),
	.d(\ctrl_opcode~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_opcode[1]~2_combout ),
	.q(ctrl_opcode_2),
	.prn(vcc));
defparam \ctrl_opcode[2] .is_wysiwyg = "true";
defparam \ctrl_opcode[2] .power_up = "low";

dffeas \ctrl_opcode[0] (
	.clk(clk),
	.d(\ctrl_opcode~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_opcode_0),
	.prn(vcc));
defparam \ctrl_opcode[0] .is_wysiwyg = "true";
defparam \ctrl_opcode[0] .power_up = "low";

dffeas ctrl_go(
	.clk(clk),
	.d(\ctrl_opcode[1]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_go1),
	.prn(vcc));
defparam ctrl_go.is_wysiwyg = "true";
defparam ctrl_go.power_up = "low";

dffeas ctrl_lock(
	.clk(clk),
	.d(\ctrl_lock~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_lock1),
	.prn(vcc));
defparam ctrl_lock.is_wysiwyg = "true";
defparam ctrl_lock.power_up = "low";

cyclonev_lcell_comb \ctrl_op_done~0 (
	.dataa(!\rmw_offset~q ),
	.datab(!\uif_ctrl_req~q ),
	.datac(!\chn_chk_active~q ),
	.datad(!av_ctrl_req),
	.datae(!\Selector5~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_op_done),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_op_done~0 .extended_lut = "off";
defparam \ctrl_op_done~0 .lut_mask = 64'h00002FAF00002FAF;
defparam \ctrl_op_done~0 .shared_arith = "off";

dffeas \mif_err_reg[4] (
	.clk(clk),
	.d(\mif_err_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mif_err_reg_4),
	.prn(vcc));
defparam \mif_err_reg[4] .is_wysiwyg = "true";
defparam \mif_err_reg[4] .power_up = "low";

dffeas \mif_err_reg[1] (
	.clk(clk),
	.d(\mif_err_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mif_err_reg_1),
	.prn(vcc));
defparam \mif_err_reg[1] .is_wysiwyg = "true";
defparam \mif_err_reg[1] .power_up = "low";

dffeas \mif_err_reg[0] (
	.clk(clk),
	.d(\mif_err_reg~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mif_err_reg_0),
	.prn(vcc));
defparam \mif_err_reg[0] .is_wysiwyg = "true";
defparam \mif_err_reg[0] .power_up = "low";

dffeas ctrl_av_go(
	.clk(clk),
	.d(\ctrl_av_go~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_av_go1),
	.prn(vcc));
defparam ctrl_av_go.is_wysiwyg = "true";
defparam ctrl_av_go.power_up = "low";

dffeas \mif_base_addr[0] (
	.clk(clk),
	.d(uif_writedata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_0),
	.prn(vcc));
defparam \mif_base_addr[0] .is_wysiwyg = "true";
defparam \mif_base_addr[0] .power_up = "low";

dffeas \mif_base_addr[1] (
	.clk(clk),
	.d(uif_writedata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_1),
	.prn(vcc));
defparam \mif_base_addr[1] .is_wysiwyg = "true";
defparam \mif_base_addr[1] .power_up = "low";

dffeas \mif_base_addr[2] (
	.clk(clk),
	.d(uif_writedata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_2),
	.prn(vcc));
defparam \mif_base_addr[2] .is_wysiwyg = "true";
defparam \mif_base_addr[2] .power_up = "low";

dffeas \mif_base_addr[3] (
	.clk(clk),
	.d(uif_writedata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_3),
	.prn(vcc));
defparam \mif_base_addr[3] .is_wysiwyg = "true";
defparam \mif_base_addr[3] .power_up = "low";

dffeas \mif_base_addr[4] (
	.clk(clk),
	.d(uif_writedata_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_4),
	.prn(vcc));
defparam \mif_base_addr[4] .is_wysiwyg = "true";
defparam \mif_base_addr[4] .power_up = "low";

dffeas \mif_base_addr[5] (
	.clk(clk),
	.d(uif_writedata_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_5),
	.prn(vcc));
defparam \mif_base_addr[5] .is_wysiwyg = "true";
defparam \mif_base_addr[5] .power_up = "low";

dffeas \mif_base_addr[6] (
	.clk(clk),
	.d(uif_writedata_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_6),
	.prn(vcc));
defparam \mif_base_addr[6] .is_wysiwyg = "true";
defparam \mif_base_addr[6] .power_up = "low";

dffeas \mif_base_addr[7] (
	.clk(clk),
	.d(uif_writedata_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_7),
	.prn(vcc));
defparam \mif_base_addr[7] .is_wysiwyg = "true";
defparam \mif_base_addr[7] .power_up = "low";

dffeas \mif_base_addr[8] (
	.clk(clk),
	.d(uif_writedata_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_8),
	.prn(vcc));
defparam \mif_base_addr[8] .is_wysiwyg = "true";
defparam \mif_base_addr[8] .power_up = "low";

dffeas \mif_base_addr[9] (
	.clk(clk),
	.d(uif_writedata_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_9),
	.prn(vcc));
defparam \mif_base_addr[9] .is_wysiwyg = "true";
defparam \mif_base_addr[9] .power_up = "low";

dffeas \mif_base_addr[10] (
	.clk(clk),
	.d(uif_writedata_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_10),
	.prn(vcc));
defparam \mif_base_addr[10] .is_wysiwyg = "true";
defparam \mif_base_addr[10] .power_up = "low";

dffeas \mif_base_addr[11] (
	.clk(clk),
	.d(uif_writedata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_11),
	.prn(vcc));
defparam \mif_base_addr[11] .is_wysiwyg = "true";
defparam \mif_base_addr[11] .power_up = "low";

dffeas \mif_base_addr[12] (
	.clk(clk),
	.d(uif_writedata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_12),
	.prn(vcc));
defparam \mif_base_addr[12] .is_wysiwyg = "true";
defparam \mif_base_addr[12] .power_up = "low";

dffeas \mif_base_addr[13] (
	.clk(clk),
	.d(uif_writedata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_13),
	.prn(vcc));
defparam \mif_base_addr[13] .is_wysiwyg = "true";
defparam \mif_base_addr[13] .power_up = "low";

dffeas \mif_base_addr[14] (
	.clk(clk),
	.d(uif_writedata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_14),
	.prn(vcc));
defparam \mif_base_addr[14] .is_wysiwyg = "true";
defparam \mif_base_addr[14] .power_up = "low";

dffeas \mif_base_addr[15] (
	.clk(clk),
	.d(uif_writedata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_15),
	.prn(vcc));
defparam \mif_base_addr[15] .is_wysiwyg = "true";
defparam \mif_base_addr[15] .power_up = "low";

dffeas \mif_base_addr[16] (
	.clk(clk),
	.d(uif_writedata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_16),
	.prn(vcc));
defparam \mif_base_addr[16] .is_wysiwyg = "true";
defparam \mif_base_addr[16] .power_up = "low";

dffeas \mif_base_addr[17] (
	.clk(clk),
	.d(uif_writedata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_17),
	.prn(vcc));
defparam \mif_base_addr[17] .is_wysiwyg = "true";
defparam \mif_base_addr[17] .power_up = "low";

dffeas \mif_base_addr[18] (
	.clk(clk),
	.d(uif_writedata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_18),
	.prn(vcc));
defparam \mif_base_addr[18] .is_wysiwyg = "true";
defparam \mif_base_addr[18] .power_up = "low";

dffeas \mif_base_addr[19] (
	.clk(clk),
	.d(uif_writedata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_19),
	.prn(vcc));
defparam \mif_base_addr[19] .is_wysiwyg = "true";
defparam \mif_base_addr[19] .power_up = "low";

dffeas \mif_base_addr[20] (
	.clk(clk),
	.d(uif_writedata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_20),
	.prn(vcc));
defparam \mif_base_addr[20] .is_wysiwyg = "true";
defparam \mif_base_addr[20] .power_up = "low";

dffeas \mif_base_addr[21] (
	.clk(clk),
	.d(uif_writedata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_21),
	.prn(vcc));
defparam \mif_base_addr[21] .is_wysiwyg = "true";
defparam \mif_base_addr[21] .power_up = "low";

dffeas \mif_base_addr[22] (
	.clk(clk),
	.d(uif_writedata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_22),
	.prn(vcc));
defparam \mif_base_addr[22] .is_wysiwyg = "true";
defparam \mif_base_addr[22] .power_up = "low";

dffeas \mif_base_addr[23] (
	.clk(clk),
	.d(uif_writedata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_23),
	.prn(vcc));
defparam \mif_base_addr[23] .is_wysiwyg = "true";
defparam \mif_base_addr[23] .power_up = "low";

dffeas \mif_base_addr[24] (
	.clk(clk),
	.d(uif_writedata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_24),
	.prn(vcc));
defparam \mif_base_addr[24] .is_wysiwyg = "true";
defparam \mif_base_addr[24] .power_up = "low";

dffeas \mif_base_addr[25] (
	.clk(clk),
	.d(uif_writedata_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_25),
	.prn(vcc));
defparam \mif_base_addr[25] .is_wysiwyg = "true";
defparam \mif_base_addr[25] .power_up = "low";

dffeas \mif_base_addr[26] (
	.clk(clk),
	.d(uif_writedata_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_26),
	.prn(vcc));
defparam \mif_base_addr[26] .is_wysiwyg = "true";
defparam \mif_base_addr[26] .power_up = "low";

dffeas \mif_base_addr[27] (
	.clk(clk),
	.d(uif_writedata_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_27),
	.prn(vcc));
defparam \mif_base_addr[27] .is_wysiwyg = "true";
defparam \mif_base_addr[27] .power_up = "low";

dffeas \mif_base_addr[28] (
	.clk(clk),
	.d(uif_writedata_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_28),
	.prn(vcc));
defparam \mif_base_addr[28] .is_wysiwyg = "true";
defparam \mif_base_addr[28] .power_up = "low";

dffeas \mif_base_addr[29] (
	.clk(clk),
	.d(uif_writedata_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_29),
	.prn(vcc));
defparam \mif_base_addr[29] .is_wysiwyg = "true";
defparam \mif_base_addr[29] .power_up = "low";

dffeas \mif_base_addr[30] (
	.clk(clk),
	.d(uif_writedata_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_30),
	.prn(vcc));
defparam \mif_base_addr[30] .is_wysiwyg = "true";
defparam \mif_base_addr[30] .power_up = "low";

dffeas \mif_base_addr[31] (
	.clk(clk),
	.d(uif_writedata_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_base_addr[31]~0_combout ),
	.q(mif_base_addr_31),
	.prn(vcc));
defparam \mif_base_addr[31] .is_wysiwyg = "true";
defparam \mif_base_addr[31] .power_up = "low";

dffeas \ctrl_wdata[1] (
	.clk(clk),
	.d(\ctrl_wdata~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_1),
	.prn(vcc));
defparam \ctrl_wdata[1] .is_wysiwyg = "true";
defparam \ctrl_wdata[1] .power_up = "low";

dffeas \ctrl_wdata[2] (
	.clk(clk),
	.d(\ctrl_wdata~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_2),
	.prn(vcc));
defparam \ctrl_wdata[2] .is_wysiwyg = "true";
defparam \ctrl_wdata[2] .power_up = "low";

dffeas \ctrl_wdata[0] (
	.clk(clk),
	.d(\ctrl_wdata~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_0),
	.prn(vcc));
defparam \ctrl_wdata[0] .is_wysiwyg = "true";
defparam \ctrl_wdata[0] .power_up = "low";

dffeas \ctrl_wdata[3] (
	.clk(clk),
	.d(\ctrl_wdata~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_3),
	.prn(vcc));
defparam \ctrl_wdata[3] .is_wysiwyg = "true";
defparam \ctrl_wdata[3] .power_up = "low";

dffeas \ctrl_addr[3] (
	.clk(clk),
	.d(\ctrl_addr~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_addr~2_combout ),
	.q(ctrl_addr_3),
	.prn(vcc));
defparam \ctrl_addr[3] .is_wysiwyg = "true";
defparam \ctrl_addr[3] .power_up = "low";

dffeas \ctrl_wdata[4] (
	.clk(clk),
	.d(\ctrl_wdata~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_4),
	.prn(vcc));
defparam \ctrl_wdata[4] .is_wysiwyg = "true";
defparam \ctrl_wdata[4] .power_up = "low";

dffeas \ctrl_wdata[5] (
	.clk(clk),
	.d(\ctrl_wdata~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_5),
	.prn(vcc));
defparam \ctrl_wdata[5] .is_wysiwyg = "true";
defparam \ctrl_wdata[5] .power_up = "low";

dffeas \ctrl_wdata[6] (
	.clk(clk),
	.d(\ctrl_wdata~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_6),
	.prn(vcc));
defparam \ctrl_wdata[6] .is_wysiwyg = "true";
defparam \ctrl_wdata[6] .power_up = "low";

dffeas \ctrl_wdata[7] (
	.clk(clk),
	.d(\ctrl_wdata~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_7),
	.prn(vcc));
defparam \ctrl_wdata[7] .is_wysiwyg = "true";
defparam \ctrl_wdata[7] .power_up = "low";

dffeas \ctrl_wdata[8] (
	.clk(clk),
	.d(\ctrl_wdata~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_8),
	.prn(vcc));
defparam \ctrl_wdata[8] .is_wysiwyg = "true";
defparam \ctrl_wdata[8] .power_up = "low";

dffeas \ctrl_wdata[9] (
	.clk(clk),
	.d(\ctrl_wdata~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_9),
	.prn(vcc));
defparam \ctrl_wdata[9] .is_wysiwyg = "true";
defparam \ctrl_wdata[9] .power_up = "low";

dffeas \ctrl_wdata[10] (
	.clk(clk),
	.d(\ctrl_wdata~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_10),
	.prn(vcc));
defparam \ctrl_wdata[10] .is_wysiwyg = "true";
defparam \ctrl_wdata[10] .power_up = "low";

dffeas \ctrl_wdata[11] (
	.clk(clk),
	.d(\ctrl_wdata~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_11),
	.prn(vcc));
defparam \ctrl_wdata[11] .is_wysiwyg = "true";
defparam \ctrl_wdata[11] .power_up = "low";

dffeas \ctrl_addr[11] (
	.clk(clk),
	.d(\ctrl_addr~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_addr~2_combout ),
	.q(ctrl_addr_11),
	.prn(vcc));
defparam \ctrl_addr[11] .is_wysiwyg = "true";
defparam \ctrl_addr[11] .power_up = "low";

dffeas \ctrl_wdata[12] (
	.clk(clk),
	.d(\ctrl_wdata~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_12),
	.prn(vcc));
defparam \ctrl_wdata[12] .is_wysiwyg = "true";
defparam \ctrl_wdata[12] .power_up = "low";

dffeas \ctrl_wdata[13] (
	.clk(clk),
	.d(\ctrl_wdata~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_13),
	.prn(vcc));
defparam \ctrl_wdata[13] .is_wysiwyg = "true";
defparam \ctrl_wdata[13] .power_up = "low";

dffeas \ctrl_wdata[14] (
	.clk(clk),
	.d(\ctrl_wdata~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_14),
	.prn(vcc));
defparam \ctrl_wdata[14] .is_wysiwyg = "true";
defparam \ctrl_wdata[14] .power_up = "low";

dffeas \ctrl_wdata[15] (
	.clk(clk),
	.d(\ctrl_wdata~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_wdata_15),
	.prn(vcc));
defparam \ctrl_wdata[15] .is_wysiwyg = "true";
defparam \ctrl_wdata[15] .power_up = "low";

dffeas mif_addr_mode(
	.clk(clk),
	.d(\mif_addr_mode~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mif_addr_mode1),
	.prn(vcc));
defparam mif_addr_mode.is_wysiwyg = "true";
defparam mif_addr_mode.power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~0 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~0 .extended_lut = "off";
defparam \ctrl_wdata~0 .lut_mask = 64'h8888888888888888;
defparam \ctrl_wdata~0 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!uif_go),
	.datad(!\ctrl_wdata~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'h0008000800080008;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_addr_offset_1),
	.datac(!uif_addr_offset_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h8080808080808080;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata[11]~3 (
	.dataa(!\always1~0_combout ),
	.datab(!\Equal3~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata[11]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata[11]~3 .extended_lut = "off";
defparam \uif_rdata[11]~3 .lut_mask = 64'h4444444444444444;
defparam \uif_rdata[11]~3 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata[2]~0 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!uif_go),
	.datad(!\ctrl_wdata~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata[2]~0 .extended_lut = "off";
defparam \uif_rdata[2]~0 .lut_mask = 64'h8808880888088808;
defparam \uif_rdata[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!Equal5),
	.datab(!uif_go),
	.datac(!\ctrl_wdata~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0101010101010101;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_strm_start~0 (
	.dataa(!uif_writedata_0),
	.datab(!\always0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_strm_start~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_strm_start~0 .extended_lut = "off";
defparam \mif_strm_start~0 .lut_mask = 64'h1111111111111111;
defparam \mif_strm_start~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_strm_start~1 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_addr_offset_1),
	.datac(!uif_addr_offset_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_strm_start~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_strm_start~1 .extended_lut = "off";
defparam \mif_strm_start~1 .lut_mask = 64'hFF40FF40FF40FF40;
defparam \mif_strm_start~1 .shared_arith = "off";

dffeas mif_strm_start(
	.clk(clk),
	.d(\mif_strm_start~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_strm_start~1_combout ),
	.q(\mif_strm_start~q ),
	.prn(vcc));
defparam mif_strm_start.is_wysiwyg = "true";
defparam mif_strm_start.power_up = "low";

cyclonev_lcell_comb \ctrl_next_state~0 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!uif_go),
	.datad(!\ctrl_wdata~0_combout ),
	.datae(!\mif_strm_start~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_next_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_next_state~0 .extended_lut = "off";
defparam \ctrl_next_state~0 .lut_mask = 64'h0C040C000C040C00;
defparam \ctrl_next_state~0 .shared_arith = "off";

cyclonev_lcell_comb \set_uif_ctrl_req~0 (
	.dataa(!Equal5),
	.datab(!\ctrl_state.CTRL_IDLE~q ),
	.datac(!uif_go),
	.datad(!\ctrl_wdata~0_combout ),
	.datae(!\ctrl_next_state~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\set_uif_ctrl_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \set_uif_ctrl_req~0 .extended_lut = "off";
defparam \set_uif_ctrl_req~0 .lut_mask = 64'h0400CCCC0400CCCC;
defparam \set_uif_ctrl_req~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_ctrl_req~0 (
	.dataa(!\uif_ctrl_req~q ),
	.datab(!ctrl_op_done),
	.datac(!\set_uif_ctrl_req~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_ctrl_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_ctrl_req~0 .extended_lut = "off";
defparam \uif_ctrl_req~0 .lut_mask = 64'h4F4F4F4F4F4F4F4F;
defparam \uif_ctrl_req~0 .shared_arith = "off";

dffeas uif_ctrl_req(
	.clk(clk),
	.d(\uif_ctrl_req~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\uif_ctrl_req~q ),
	.prn(vcc));
defparam uif_ctrl_req.is_wysiwyg = "true";
defparam uif_ctrl_req.power_up = "low";

cyclonev_lcell_comb \chn_chk_active~0 (
	.dataa(!\chn_chk_active~q ),
	.datab(!\Selector5~1_combout ),
	.datac(!\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\chn_chk_active~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \chn_chk_active~0 .extended_lut = "off";
defparam \chn_chk_active~0 .lut_mask = 64'h4F4F4F4F4F4F4F4F;
defparam \chn_chk_active~0 .shared_arith = "off";

dffeas chn_chk_active(
	.clk(clk),
	.d(\chn_chk_active~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\chn_chk_active~q ),
	.prn(vcc));
defparam chn_chk_active.is_wysiwyg = "true";
defparam chn_chk_active.power_up = "low";

cyclonev_lcell_comb \always3~0 (
	.dataa(!\rmw_offset~q ),
	.datab(!\chn_chk_active~q ),
	.datac(!av_ctrl_req),
	.datad(!waitrequest_to_ctrl),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~0 .extended_lut = "off";
defparam \always3~0 .lut_mask = 64'h3B003B003B003B00;
defparam \always3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!av_ctrl_req),
	.datab(!\ctrl_state.CTRL_WF_B~q ),
	.datac(!av_done),
	.datad(!\ctrl_state.CTRL_WF_AV~q ),
	.datae(!\always3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h00A033B300A033B3;
defparam \Selector8~0 .shared_arith = "off";

dffeas \ctrl_state.CTRL_WF_AV (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_WF_AV~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_WF_AV .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_WF_AV .power_up = "low";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!Equal5),
	.datab(!\ctrl_state.CTRL_IDLE~q ),
	.datac(!uif_go),
	.datad(!\ctrl_wdata~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h0400040004000400;
defparam \Selector10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~1 (
	.dataa(!av_ctrl_req),
	.datab(!av_done),
	.datac(!\ctrl_state.CTRL_WF_AV~q ),
	.datad(!\Selector10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~1 .extended_lut = "off";
defparam \Selector10~1 .lut_mask = 64'h04FF04FF04FF04FF;
defparam \Selector10~1 .shared_arith = "off";

dffeas \ctrl_state.CTRL_CHK_ADDR (
	.clk(clk),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_CHK_ADDR~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_CHK_ADDR .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_CHK_ADDR .power_up = "low";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!\rmw_offset~q ),
	.datab(!\ctrl_state.CTRL_CHK_ADDR~q ),
	.datac(!\ctrl_state.CTRL_RMW~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \Selector6~0 .shared_arith = "off";

dffeas \ctrl_state.CTRL_MIF_WR (
	.clk(clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_MIF_WR~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_MIF_WR .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_MIF_WR .power_up = "low";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!\rmw_offset~q ),
	.datab(!\ctrl_state.CTRL_IDLE~q ),
	.datac(!\ctrl_state.CTRL_CHK_ADDR~q ),
	.datad(!\ctrl_next_state~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector9~0 .shared_arith = "off";

dffeas \ctrl_state.CTRL_MIF_RD (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_MIF_RD~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_MIF_RD .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_MIF_RD .power_up = "low";

dffeas \ctrl_state.CTRL_CHK_CHN (
	.clk(clk),
	.d(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_CHK_CHN~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_CHK_CHN .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_CHK_CHN .power_up = "low";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!\uif_ctrl_req~q ),
	.datab(!\chn_chk_active~q ),
	.datac(!av_ctrl_req),
	.datad(!waitrequest_to_ctrl),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h7F007F007F007F00;
defparam \Selector7~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~1 (
	.dataa(!\ctrl_state.CTRL_WF_B~q ),
	.datab(!\ctrl_state.CTRL_MIF_WR~q ),
	.datac(!\ctrl_state.CTRL_MIF_RD~q ),
	.datad(!\ctrl_state.CTRL_CHK_CHN~q ),
	.datae(!\Selector7~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~1 .extended_lut = "off";
defparam \Selector7~1 .lut_mask = 64'h7FFF3FFF7FFF3FFF;
defparam \Selector7~1 .shared_arith = "off";

dffeas \ctrl_state.CTRL_WF_B (
	.clk(clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_WF_B~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_WF_B .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_WF_B .power_up = "low";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!waitrequest_to_ctrl),
	.datab(!\ctrl_state.CTRL_WF_B~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'h2222222222222222;
defparam \Selector5~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_next_state.CTRL_RMW~0 (
	.dataa(!\rmw_offset~q ),
	.datab(!\uif_ctrl_req~q ),
	.datac(!av_ctrl_req),
	.datad(!\Selector5~1_combout ),
	.datae(!\always3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_next_state.CTRL_RMW~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_next_state.CTRL_RMW~0 .extended_lut = "off";
defparam \ctrl_next_state.CTRL_RMW~0 .lut_mask = 64'h0015000000150000;
defparam \ctrl_next_state.CTRL_RMW~0 .shared_arith = "off";

dffeas \ctrl_state.CTRL_RMW (
	.clk(clk),
	.d(\ctrl_next_state.CTRL_RMW~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_RMW~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_RMW .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_RMW .power_up = "low";

dffeas av_ctrl_req_dly(
	.clk(clk),
	.d(av_ctrl_req),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ctrl_req_dly~q ),
	.prn(vcc));
defparam av_ctrl_req_dly.is_wysiwyg = "true";
defparam av_ctrl_req_dly.power_up = "low";

cyclonev_lcell_comb \always9~0 (
	.dataa(!Equal5),
	.datab(!uif_ctrl_0),
	.datac(!uif_ctrl_1),
	.datad(!av_ctrl_req),
	.datae(!uif_go),
	.dataf(!\av_ctrl_req_dly~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~0 .extended_lut = "off";
defparam \always9~0 .lut_mask = 64'h00FF10FF00001010;
defparam \always9~0 .shared_arith = "off";

cyclonev_lcell_comb \mux_mif_addr[4]~0 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_4),
	.datad(!av_mif_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_mif_addr[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_mif_addr[4]~0 .extended_lut = "off";
defparam \mux_mif_addr[4]~0 .lut_mask = 64'h078F078F078F078F;
defparam \mux_mif_addr[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \mux_mif_addr[5]~1 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_5),
	.datad(!av_mif_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_mif_addr[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_mif_addr[5]~1 .extended_lut = "off";
defparam \mux_mif_addr[5]~1 .lut_mask = 64'h078F078F078F078F;
defparam \mux_mif_addr[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \mux_mif_addr[2]~2 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_addr_offset_2),
	.datac(!uif_ctrl_1),
	.datad(!av_mif_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_mif_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_mif_addr[2]~2 .extended_lut = "off";
defparam \mux_mif_addr[2]~2 .lut_mask = 64'h13B313B313B313B3;
defparam \mux_mif_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \mux_mif_addr[1]~3 (
	.dataa(!uif_addr_offset_1),
	.datab(!uif_ctrl_0),
	.datac(!uif_ctrl_1),
	.datad(!av_mif_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_mif_addr[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_mif_addr[1]~3 .extended_lut = "off";
defparam \mux_mif_addr[1]~3 .lut_mask = 64'h15D515D515D515D5;
defparam \mux_mif_addr[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \mux_mif_addr[0]~4 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_ctrl_0),
	.datac(!uif_ctrl_1),
	.datad(!av_mif_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_mif_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_mif_addr[0]~4 .extended_lut = "off";
defparam \mux_mif_addr[0]~4 .lut_mask = 64'h15D515D515D515D5;
defparam \mux_mif_addr[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \mux_mif_addr[3]~5 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_3),
	.datad(!av_mif_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_mif_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_mif_addr[3]~5 .extended_lut = "off";
defparam \mux_mif_addr[3]~5 .lut_mask = 64'h078F078F078F078F;
defparam \mux_mif_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~0 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_8),
	.datad(!uif_addr_offset_9),
	.datae(!uif_addr_offset_11),
	.dataf(!av_mif_addr_8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'hF888888870000000;
defparam \Equal14~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~1 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_10),
	.datad(!av_mif_addr_9),
	.datae(!av_mif_addr_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~1 .extended_lut = "off";
defparam \Equal14~1 .lut_mask = 64'hF8707070F8707070;
defparam \Equal14~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~2 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_6),
	.datad(!uif_addr_offset_7),
	.datae(!av_mif_addr_7),
	.dataf(!av_mif_addr_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~2 .extended_lut = "off";
defparam \Equal14~2 .lut_mask = 64'hF888700070007000;
defparam \Equal14~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~3 (
	.dataa(!\mux_mif_addr[0]~4_combout ),
	.datab(!\mux_mif_addr[3]~5_combout ),
	.datac(!\Equal14~0_combout ),
	.datad(!\Equal14~1_combout ),
	.datae(!\Equal14~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~3 .extended_lut = "off";
defparam \Equal14~3 .lut_mask = 64'h0000000800000008;
defparam \Equal14~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal22~0 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_4),
	.datad(!uif_addr_offset_5),
	.datae(!av_mif_addr_4),
	.dataf(!av_mif_addr_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~0 .extended_lut = "off";
defparam \Equal22~0 .lut_mask = 64'hF888700070007000;
defparam \Equal22~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal22~1 (
	.dataa(!uif_addr_offset_1),
	.datab(!uif_ctrl_0),
	.datac(!uif_addr_offset_2),
	.datad(!uif_ctrl_1),
	.datae(!av_mif_addr_2),
	.dataf(!av_mif_addr_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~1 .extended_lut = "off";
defparam \Equal22~1 .lut_mask = 64'h010501050105CD05;
defparam \Equal22~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~0 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_ctrl_0),
	.datac(!uif_ctrl_1),
	.datad(!uif_addr_offset_3),
	.datae(!av_mif_addr_0),
	.dataf(!av_mif_addr_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~0 .extended_lut = "off";
defparam \Equal17~0 .lut_mask = 64'h001500150015C0D5;
defparam \Equal17~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~1 (
	.dataa(!\Equal14~0_combout ),
	.datab(!\Equal14~1_combout ),
	.datac(!\Equal14~2_combout ),
	.datad(!\Equal22~0_combout ),
	.datae(!\Equal22~1_combout ),
	.dataf(!\Equal17~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~1 .extended_lut = "off";
defparam \Equal17~1 .lut_mask = 64'h0000000000000001;
defparam \Equal17~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~1 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~1 .extended_lut = "off";
defparam \ctrl_wdata~1 .lut_mask = 64'hFFFF7DFF00000000;
defparam \ctrl_wdata~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~4 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~4 .extended_lut = "off";
defparam \Equal14~4 .lut_mask = 64'h8080808080808080;
defparam \Equal14~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~5 (
	.dataa(!\mux_mif_addr[3]~5_combout ),
	.datab(!\Equal14~0_combout ),
	.datac(!\Equal14~1_combout ),
	.datad(!\Equal14~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~5 .extended_lut = "off";
defparam \Equal14~5 .lut_mask = 64'h0002000200020002;
defparam \Equal14~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~0 (
	.dataa(!\Equal14~4_combout ),
	.datab(!\mux_mif_addr[1]~3_combout ),
	.datac(!\mux_mif_addr[0]~4_combout ),
	.datad(!\Equal14~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~0 .extended_lut = "off";
defparam \Equal15~0 .lut_mask = 64'h0004000400040004;
defparam \Equal15~0 .shared_arith = "off";

cyclonev_lcell_comb \mux_mif_addr[6]~6 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_6),
	.datad(!av_mif_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_mif_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_mif_addr[6]~6 .extended_lut = "off";
defparam \mux_mif_addr[6]~6 .lut_mask = 64'h078F078F078F078F;
defparam \mux_mif_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal23~0 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_addr_offset_3),
	.datad(!uif_addr_offset_7),
	.datae(!av_mif_addr_3),
	.dataf(!av_mif_addr_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~0 .extended_lut = "off";
defparam \Equal23~0 .lut_mask = 64'h000700070007888F;
defparam \Equal23~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal23~1 (
	.dataa(!\mux_mif_addr[1]~3_combout ),
	.datab(!\mux_mif_addr[0]~4_combout ),
	.datac(!\mux_mif_addr[6]~6_combout ),
	.datad(!\Equal14~0_combout ),
	.datae(!\Equal14~1_combout ),
	.dataf(!\Equal23~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~1 .extended_lut = "off";
defparam \Equal23~1 .lut_mask = 64'h0000000000000004;
defparam \Equal23~1 .shared_arith = "off";

cyclonev_lcell_comb \WideNor1~0 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal23~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~0 .extended_lut = "off";
defparam \WideNor1~0 .lut_mask = 64'h000040E8404040E8;
defparam \WideNor1~0 .shared_arith = "off";

cyclonev_lcell_comb \rmw_offset~0 (
	.dataa(!\rmw_offset~q ),
	.datab(!\ctrl_state.CTRL_RMW~q ),
	.datac(!\always9~0_combout ),
	.datad(!\ctrl_wdata~1_combout ),
	.datae(!\Equal15~0_combout ),
	.dataf(!\WideNor1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rmw_offset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rmw_offset~0 .extended_lut = "off";
defparam \rmw_offset~0 .lut_mask = 64'h4C404C4C4C4C4C4C;
defparam \rmw_offset~0 .shared_arith = "off";

dffeas rmw_offset(
	.clk(clk),
	.d(\rmw_offset~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rmw_offset~q ),
	.prn(vcc));
defparam rmw_offset.is_wysiwyg = "true";
defparam rmw_offset.power_up = "low";

cyclonev_lcell_comb \ctrl_next_state~1 (
	.dataa(!\rmw_offset~q ),
	.datab(!\uif_ctrl_req~q ),
	.datac(!\chn_chk_active~q ),
	.datad(!av_ctrl_req),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_next_state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_next_state~1 .extended_lut = "off";
defparam \ctrl_next_state~1 .lut_mask = 64'h2000200020002000;
defparam \ctrl_next_state~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~2 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!\ctrl_state.CTRL_IDLE~q ),
	.datad(!uif_go),
	.datae(!\ctrl_wdata~0_combout ),
	.dataf(!\mif_strm_start~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~2 .extended_lut = "off";
defparam \Selector5~2 .lut_mask = 64'hF010F0B0F0100000;
defparam \Selector5~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~3 (
	.dataa(!\ctrl_next_state~1_combout ),
	.datab(!\Selector5~1_combout ),
	.datac(!av_done),
	.datad(!\ctrl_state.CTRL_WF_AV~q ),
	.datae(!\Selector5~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~3 .extended_lut = "off";
defparam \Selector5~3 .lut_mask = 64'hEEE00000EEE00000;
defparam \Selector5~3 .shared_arith = "off";

dffeas \ctrl_state.CTRL_IDLE (
	.clk(clk),
	.d(\Selector5~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CTRL_IDLE~q ),
	.prn(vcc));
defparam \ctrl_state.CTRL_IDLE .is_wysiwyg = "true";
defparam \ctrl_state.CTRL_IDLE .power_up = "low";

cyclonev_lcell_comb \ctrl_next_state.CTRL_CHK_CHN~0 (
	.dataa(!\ctrl_state.CTRL_IDLE~q ),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!\mif_strm_start~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_next_state.CTRL_CHK_CHN~0 .extended_lut = "off";
defparam \ctrl_next_state.CTRL_CHK_CHN~0 .lut_mask = 64'h0202020202020202;
defparam \ctrl_next_state.CTRL_CHK_CHN~0 .shared_arith = "off";

cyclonev_lcell_comb \always6~0 (
	.dataa(!av_ctrl_req),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!\av_ctrl_req_dly~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \always6~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr[1]~0 (
	.dataa(!av_ctrl_req),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.datad(!\av_ctrl_req_dly~q ),
	.datae(!\set_uif_ctrl_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr[1]~0 .extended_lut = "off";
defparam \ctrl_addr[1]~0 .lut_mask = 64'h1F0FDFCF1F0FDFCF;
defparam \ctrl_addr[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~12 (
	.dataa(!uif_addr_offset_2),
	.datab(!uif_addr_offset_0),
	.datac(!mif_err_reg_0),
	.datad(!\always1~0_combout ),
	.datae(!uif_addr_offset_1),
	.dataf(!ctrl_rdata[0]),
	.datag(!mif_base_addr_0),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~12 .extended_lut = "on";
defparam \uif_rdata~12 .lut_mask = 64'h00080008FF08FF08;
defparam \uif_rdata~12 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~8 (
	.dataa(!uif_addr_offset_2),
	.datab(!uif_addr_offset_0),
	.datac(!mif_err_reg_1),
	.datad(!ctrl_rdata[1]),
	.datae(!uif_addr_offset_1),
	.dataf(!\always1~0_combout ),
	.datag(!mif_base_addr_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~8 .extended_lut = "on";
defparam \uif_rdata~8 .lut_mask = 64'h00FF00FF08080808;
defparam \uif_rdata~8 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~1 (
	.dataa(!mif_base_addr_2),
	.datab(!\always1~0_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!ctrl_rdata[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~1 .extended_lut = "off";
defparam \uif_rdata~1 .lut_mask = 64'h01CD01CD01CD01CD;
defparam \uif_rdata~1 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~2 (
	.dataa(!mif_base_addr_3),
	.datab(!\always1~0_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!ctrl_rdata[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~2 .extended_lut = "off";
defparam \uif_rdata~2 .lut_mask = 64'h01CD01CD01CD01CD;
defparam \uif_rdata~2 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~4 (
	.dataa(!uif_addr_offset_2),
	.datab(!uif_addr_offset_0),
	.datac(!mif_err_reg_4),
	.datad(!ctrl_rdata[4]),
	.datae(!uif_addr_offset_1),
	.dataf(!\always1~0_combout ),
	.datag(!mif_base_addr_4),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~4 .extended_lut = "on";
defparam \uif_rdata~4 .lut_mask = 64'h00FF00FF08080808;
defparam \uif_rdata~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!uif_addr_offset_7),
	.datab(!uif_addr_offset_8),
	.datac(!uif_addr_offset_9),
	.datad(!uif_addr_offset_10),
	.datae(!uif_addr_offset_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8000000080000000;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!uif_addr_offset_2),
	.datab(!uif_addr_offset_3),
	.datac(!uif_addr_offset_4),
	.datad(!uif_addr_offset_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h8000800080008000;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb uif_addr_err_d(
	.dataa(!uif_addr_offset_0),
	.datab(!uif_addr_offset_1),
	.datac(!uif_addr_offset_6),
	.datad(!\ctrl_wdata~0_combout ),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\LessThan0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_addr_err_d~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam uif_addr_err_d.extended_lut = "off";
defparam uif_addr_err_d.lut_mask = 64'h00FF00FF00FF001F;
defparam uif_addr_err_d.shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode~0 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode~0 .extended_lut = "off";
defparam \ctrl_opcode~0 .lut_mask = 64'h1111111111111111;
defparam \ctrl_opcode~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode~1 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!\Selector6~0_combout ),
	.datad(!\Selector9~0_combout ),
	.datae(!\ctrl_opcode~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode~1 .extended_lut = "off";
defparam \ctrl_opcode~1 .lut_mask = 64'h00440F4F00440F4F;
defparam \ctrl_opcode~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode[1]~2 (
	.dataa(!\Selector6~0_combout ),
	.datab(!\Selector9~0_combout ),
	.datac(!\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode[1]~2 .extended_lut = "off";
defparam \ctrl_opcode[1]~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ctrl_opcode[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode~3 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!\Selector6~0_combout ),
	.datad(!\Selector9~0_combout ),
	.datae(!\ctrl_opcode~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode~3 .extended_lut = "off";
defparam \ctrl_opcode~3 .lut_mask = 64'h00000F8F00000F8F;
defparam \ctrl_opcode~3 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode~4 (
	.dataa(!\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.datab(!\ctrl_opcode~0_combout ),
	.datac(!uif_mode_1),
	.datad(!\Selector6~0_combout ),
	.datae(!\Selector9~0_combout ),
	.dataf(!uif_mode_0),
	.datag(!ctrl_opcode_0),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode~4 .extended_lut = "on";
defparam \ctrl_opcode~4 .lut_mask = 64'h0ACC30C00ACC00CC;
defparam \ctrl_opcode~4 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lock~0 (
	.dataa(!\rmw_offset~q ),
	.datab(!av_addr_burst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_lock~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lock~0 .extended_lut = "off";
defparam \ctrl_lock~0 .lut_mask = 64'h7777777777777777;
defparam \ctrl_lock~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_clr_error~0 (
	.dataa(!uif_writedata_2),
	.datab(!\always0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_clr_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_clr_error~0 .extended_lut = "off";
defparam \mif_clr_error~0 .lut_mask = 64'h1111111111111111;
defparam \mif_clr_error~0 .shared_arith = "off";

dffeas mif_clr_error(
	.clk(clk),
	.d(\mif_clr_error~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mif_strm_start~1_combout ),
	.q(\mif_clr_error~q ),
	.prn(vcc));
defparam mif_clr_error.is_wysiwyg = "true";
defparam mif_clr_error.power_up = "low";

cyclonev_lcell_comb \channel_id~2 (
	.dataa(!\ctrl_state.CTRL_IDLE~q ),
	.datab(!ctrl_rdata[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\channel_id~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \channel_id~2 .extended_lut = "off";
defparam \channel_id~2 .lut_mask = 64'h1111111111111111;
defparam \channel_id~2 .shared_arith = "off";

cyclonev_lcell_comb \always7~0 (
	.dataa(!ctrl_opcode_1),
	.datab(!ctrl_opcode_2),
	.datac(!ctrl_opcode_0),
	.datad(!waitrequest_to_ctrl),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always7~0 .extended_lut = "off";
defparam \always7~0 .lut_mask = 64'h8000800080008000;
defparam \always7~0 .shared_arith = "off";

cyclonev_lcell_comb \channel_id[0]~1 (
	.dataa(!\chn_chk_active~q ),
	.datab(!\ctrl_state.CTRL_IDLE~q ),
	.datac(!\always7~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\channel_id[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \channel_id[0]~1 .extended_lut = "off";
defparam \channel_id[0]~1 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \channel_id[0]~1 .shared_arith = "off";

dffeas \channel_id[0] (
	.clk(clk),
	.d(\channel_id~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_id[0]~1_combout ),
	.q(\channel_id[0]~q ),
	.prn(vcc));
defparam \channel_id[0] .is_wysiwyg = "true";
defparam \channel_id[0] .power_up = "low";

cyclonev_lcell_comb \channel_id~0 (
	.dataa(!\ctrl_state.CTRL_IDLE~q ),
	.datab(!ctrl_rdata[1]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\channel_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \channel_id~0 .extended_lut = "off";
defparam \channel_id~0 .lut_mask = 64'h1111111111111111;
defparam \channel_id~0 .shared_arith = "off";

dffeas \channel_id[1] (
	.clk(clk),
	.d(\channel_id~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_id[0]~1_combout ),
	.q(\channel_id[1]~q ),
	.prn(vcc));
defparam \channel_id[1] .is_wysiwyg = "true";
defparam \channel_id[1] .power_up = "low";

cyclonev_lcell_comb \channel_id~3 (
	.dataa(!\ctrl_state.CTRL_IDLE~q ),
	.datab(!ctrl_rdata[3]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\channel_id~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \channel_id~3 .extended_lut = "off";
defparam \channel_id~3 .lut_mask = 64'h1111111111111111;
defparam \channel_id~3 .shared_arith = "off";

dffeas \channel_id[3] (
	.clk(clk),
	.d(\channel_id~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_id[0]~1_combout ),
	.q(\channel_id[3]~q ),
	.prn(vcc));
defparam \channel_id[3] .is_wysiwyg = "true";
defparam \channel_id[3] .power_up = "low";

cyclonev_lcell_comb \channel_id~4 (
	.dataa(!\ctrl_state.CTRL_IDLE~q ),
	.datab(!ctrl_rdata[2]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\channel_id~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \channel_id~4 .extended_lut = "off";
defparam \channel_id~4 .lut_mask = 64'h1111111111111111;
defparam \channel_id~4 .shared_arith = "off";

dffeas \channel_id[2] (
	.clk(clk),
	.d(\channel_id~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_id[0]~1_combout ),
	.q(\channel_id[2]~q ),
	.prn(vcc));
defparam \channel_id[2] .is_wysiwyg = "true";
defparam \channel_id[2] .power_up = "low";

cyclonev_lcell_comb \av_chn_mismatch~0 (
	.dataa(!av_mif_type_0),
	.datab(!\channel_id[1]~q ),
	.datac(!\channel_id[0]~q ),
	.datad(!\channel_id[3]~q ),
	.datae(!\channel_id[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_chn_mismatch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_chn_mismatch~0 .extended_lut = "off";
defparam \av_chn_mismatch~0 .lut_mask = 64'hFDFDA8FDFDFDA8FD;
defparam \av_chn_mismatch~0 .shared_arith = "off";

cyclonev_lcell_comb \av_chn_mismatch~1 (
	.dataa(!\channel_id[0]~q ),
	.datab(!\channel_id[1]~q ),
	.datac(!av_mif_type_0),
	.datad(!av_mif_type_valid),
	.datae(!av_mif_type_1),
	.dataf(!\av_chn_mismatch~q ),
	.datag(!\av_chn_mismatch~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_chn_mismatch~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_chn_mismatch~1 .extended_lut = "on";
defparam \av_chn_mismatch~1 .lut_mask = 64'h000F00DB00FF00FF;
defparam \av_chn_mismatch~1 .shared_arith = "off";

dffeas av_chn_mismatch(
	.clk(clk),
	.d(\av_chn_mismatch~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_chn_mismatch~q ),
	.prn(vcc));
defparam av_chn_mismatch.is_wysiwyg = "true";
defparam av_chn_mismatch.power_up = "low";

cyclonev_lcell_comb \mif_err_reg~0 (
	.dataa(!uif_addr_err1),
	.datab(!mif_err_reg_4),
	.datac(!\uif_addr_err_d~combout ),
	.datad(!\mif_clr_error~q ),
	.datae(!\av_chn_mismatch~q ),
	.dataf(!av_opcode_err),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_err_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_err_reg~0 .extended_lut = "off";
defparam \mif_err_reg~0 .lut_mask = 64'h3300F70033003300;
defparam \mif_err_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_err_reg~1 (
	.dataa(!uif_addr_err1),
	.datab(!mif_err_reg_1),
	.datac(!\uif_addr_err_d~combout ),
	.datad(!\mif_clr_error~q ),
	.datae(!av_opcode_err),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_err_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_err_reg~1 .extended_lut = "off";
defparam \mif_err_reg~1 .lut_mask = 64'h3300F7003300F700;
defparam \mif_err_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \mif_err_reg~2 (
	.dataa(!uif_addr_err1),
	.datab(!mif_err_reg_0),
	.datac(!\uif_addr_err_d~combout ),
	.datad(!\mif_clr_error~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_err_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_err_reg~2 .extended_lut = "off";
defparam \mif_err_reg~2 .lut_mask = 64'h3B003B003B003B00;
defparam \mif_err_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_av_go~0 (
	.dataa(!\chn_chk_active~q ),
	.datab(!\Selector5~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_av_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_av_go~0 .extended_lut = "off";
defparam \ctrl_av_go~0 .lut_mask = 64'h1111111111111111;
defparam \ctrl_av_go~0 .shared_arith = "off";

cyclonev_lcell_comb \mif_base_addr[31]~0 (
	.dataa(!\Equal3~0_combout ),
	.datab(!\always0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_base_addr[31]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_base_addr[31]~0 .extended_lut = "off";
defparam \mif_base_addr[31]~0 .lut_mask = 64'h1111111111111111;
defparam \mif_base_addr[31]~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr16~0 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr16~0 .extended_lut = "off";
defparam \WideOr16~0 .lut_mask = 64'hFFFF3FDF00000000;
defparam \WideOr16~0 .shared_arith = "off";

dffeas \saved_read_data[1] (
	.clk(clk),
	.d(ctrl_rdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[1]~q ),
	.prn(vcc));
defparam \saved_read_data[1] .is_wysiwyg = "true";
defparam \saved_read_data[1] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~2 (
	.dataa(!uif_writedata_1),
	.datab(!uif_ctrl_0),
	.datac(!uif_ctrl_1),
	.datad(!\WideOr16~0_combout ),
	.datae(!\saved_read_data[1]~q ),
	.dataf(!mif_rec_data_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~2 .extended_lut = "off";
defparam \ctrl_wdata~2 .lut_mask = 64'h0515F51505D5F5D5;
defparam \ctrl_wdata~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal23~2 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\Equal23~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~2 .extended_lut = "off";
defparam \Equal23~2 .lut_mask = 64'h0040004000400040;
defparam \Equal23~2 .shared_arith = "off";

dffeas \saved_read_data[2] (
	.clk(clk),
	.d(ctrl_rdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[2]~q ),
	.prn(vcc));
defparam \saved_read_data[2] .is_wysiwyg = "true";
defparam \saved_read_data[2] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~3 (
	.dataa(!uif_writedata_2),
	.datab(!uif_ctrl_0),
	.datac(!uif_ctrl_1),
	.datad(!mif_rec_data_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~3 .extended_lut = "off";
defparam \ctrl_wdata~3 .lut_mask = 64'h11D111D111D111D1;
defparam \ctrl_wdata~3 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~4 (
	.dataa(!uif_writedata_2),
	.datab(!uif_ctrl_1),
	.datac(!\Equal23~2_combout ),
	.datad(!\WideOr16~0_combout ),
	.datae(!\saved_read_data[2]~q ),
	.dataf(!\ctrl_wdata~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~4 .extended_lut = "off";
defparam \ctrl_wdata~4 .lut_mask = 64'h1111DD1D11F1DDFD;
defparam \ctrl_wdata~4 .shared_arith = "off";

dffeas \saved_read_data[0] (
	.clk(clk),
	.d(ctrl_rdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[0]~q ),
	.prn(vcc));
defparam \saved_read_data[0] .is_wysiwyg = "true";
defparam \saved_read_data[0] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~5 (
	.dataa(!uif_writedata_0),
	.datab(!uif_ctrl_0),
	.datac(!uif_ctrl_1),
	.datad(!\saved_read_data[0]~q ),
	.datae(!\WideOr16~0_combout ),
	.dataf(!mif_rec_data_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~5 .extended_lut = "off";
defparam \ctrl_wdata~5 .lut_mask = 64'h05F5151505F5D5D5;
defparam \ctrl_wdata~5 .shared_arith = "off";

dffeas \saved_read_data[3] (
	.clk(clk),
	.d(ctrl_rdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[3]~q ),
	.prn(vcc));
defparam \saved_read_data[3] .is_wysiwyg = "true";
defparam \saved_read_data[3] .power_up = "low";

cyclonev_lcell_comb \WideOr14~0 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr14~0 .extended_lut = "off";
defparam \WideOr14~0 .lut_mask = 64'hFFFF7DDF00000000;
defparam \WideOr14~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~6 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_writedata_3),
	.datac(!uif_ctrl_1),
	.datad(!\saved_read_data[3]~q ),
	.datae(!\WideOr14~0_combout ),
	.dataf(!mif_rec_data_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~6 .extended_lut = "off";
defparam \ctrl_wdata~6 .lut_mask = 64'h03F3131303F3B3B3;
defparam \ctrl_wdata~6 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~1 (
	.dataa(!uif_addr_offset_3),
	.datab(!\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.datac(!av_mif_addr_3),
	.datad(!\always6~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~1 .extended_lut = "off";
defparam \ctrl_addr~1 .lut_mask = 64'h3F773F773F773F77;
defparam \ctrl_addr~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~2 (
	.dataa(!\ctrl_wdata~0_combout ),
	.datab(!\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.datac(!\set_uif_ctrl_req~0_combout ),
	.datad(!\always6~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~2 .extended_lut = "off";
defparam \ctrl_addr~2 .lut_mask = 64'hFF3BFF3BFF3BFF3B;
defparam \ctrl_addr~2 .shared_arith = "off";

dffeas \saved_read_data[4] (
	.clk(clk),
	.d(ctrl_rdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[4]~q ),
	.prn(vcc));
defparam \saved_read_data[4] .is_wysiwyg = "true";
defparam \saved_read_data[4] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~7 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_writedata_4),
	.datad(!\WideOr14~0_combout ),
	.datae(!\saved_read_data[4]~q ),
	.dataf(!mif_rec_data_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~7 .extended_lut = "off";
defparam \ctrl_wdata~7 .lut_mask = 64'h0307CF07038FCF8F;
defparam \ctrl_wdata~7 .shared_arith = "off";

cyclonev_lcell_comb WideOr14(
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr14~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr14.extended_lut = "off";
defparam WideOr14.lut_mask = 64'hFFFF7D9F00000000;
defparam WideOr14.shared_arith = "off";

dffeas \saved_read_data[5] (
	.clk(clk),
	.d(ctrl_rdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[5]~q ),
	.prn(vcc));
defparam \saved_read_data[5] .is_wysiwyg = "true";
defparam \saved_read_data[5] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~8 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_writedata_5),
	.datad(!\WideOr14~combout ),
	.datae(!\saved_read_data[5]~q ),
	.dataf(!mif_rec_data_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~8 .extended_lut = "off";
defparam \ctrl_wdata~8 .lut_mask = 64'h0307CF07038FCF8F;
defparam \ctrl_wdata~8 .shared_arith = "off";

dffeas \saved_read_data[6] (
	.clk(clk),
	.d(ctrl_rdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[6]~q ),
	.prn(vcc));
defparam \saved_read_data[6] .is_wysiwyg = "true";
defparam \saved_read_data[6] .power_up = "low";

cyclonev_lcell_comb \Equal20~0 (
	.dataa(!uif_addr_offset_4),
	.datab(!uif_addr_offset_5),
	.datac(!\ctrl_wdata~0_combout ),
	.datad(!av_mif_addr_4),
	.datae(!av_mif_addr_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~0 .extended_lut = "off";
defparam \Equal20~0 .lut_mask = 64'h20202F2020202F20;
defparam \Equal20~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata[6]~9 (
	.dataa(!uif_ctrl_1),
	.datab(!\mux_mif_addr[2]~2_combout ),
	.datac(!\mux_mif_addr[1]~3_combout ),
	.datad(!\Equal14~3_combout ),
	.datae(!\Equal17~1_combout ),
	.dataf(!\Equal20~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata[6]~9 .extended_lut = "off";
defparam \ctrl_wdata[6]~9 .lut_mask = 64'h0000AAAA0028AAAA;
defparam \ctrl_wdata[6]~9 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~10 (
	.dataa(!uif_writedata_6),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!\saved_read_data[6]~q ),
	.datad(!\ctrl_wdata[6]~9_combout ),
	.datae(!mif_rec_data_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~10 .extended_lut = "off";
defparam \ctrl_wdata~10 .lut_mask = 64'h440F770F440F770F;
defparam \ctrl_wdata~10 .shared_arith = "off";

dffeas \saved_read_data[7] (
	.clk(clk),
	.d(ctrl_rdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[7]~q ),
	.prn(vcc));
defparam \saved_read_data[7] .is_wysiwyg = "true";
defparam \saved_read_data[7] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~11 (
	.dataa(!uif_writedata_7),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!\ctrl_wdata[6]~9_combout ),
	.datad(!\saved_read_data[7]~q ),
	.datae(!mif_rec_data_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~11 .extended_lut = "off";
defparam \ctrl_wdata~11 .lut_mask = 64'h404F707F404F707F;
defparam \ctrl_wdata~11 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~12 (
	.dataa(!\mux_mif_addr[2]~2_combout ),
	.datab(!\mux_mif_addr[1]~3_combout ),
	.datac(!\Equal14~3_combout ),
	.datad(!\Equal17~1_combout ),
	.datae(!\Equal20~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~12 .extended_lut = "off";
defparam \ctrl_wdata~12 .lut_mask = 64'hFF00F900FF00F900;
defparam \ctrl_wdata~12 .shared_arith = "off";

dffeas \saved_read_data[8] (
	.clk(clk),
	.d(ctrl_rdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[8]~q ),
	.prn(vcc));
defparam \saved_read_data[8] .is_wysiwyg = "true";
defparam \saved_read_data[8] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~13 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_writedata_8),
	.datad(!mif_rec_data_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~13 .extended_lut = "off";
defparam \ctrl_wdata~13 .lut_mask = 64'h058D058D058D058D;
defparam \ctrl_wdata~13 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~14 (
	.dataa(!uif_ctrl_1),
	.datab(!uif_writedata_8),
	.datac(!\Equal15~0_combout ),
	.datad(!\ctrl_wdata~12_combout ),
	.datae(!\saved_read_data[8]~q ),
	.dataf(!\ctrl_wdata~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~14 .extended_lut = "off";
defparam \ctrl_wdata~14 .lut_mask = 64'h1111BB1B11F1BBFB;
defparam \ctrl_wdata~14 .shared_arith = "off";

dffeas \saved_read_data[9] (
	.clk(clk),
	.d(ctrl_rdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[9]~q ),
	.prn(vcc));
defparam \saved_read_data[9] .is_wysiwyg = "true";
defparam \saved_read_data[9] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~15 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_writedata_9),
	.datad(!mif_rec_data_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~15 .extended_lut = "off";
defparam \ctrl_wdata~15 .lut_mask = 64'h058D058D058D058D;
defparam \ctrl_wdata~15 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~16 (
	.dataa(!uif_ctrl_1),
	.datab(!uif_writedata_9),
	.datac(!\ctrl_wdata~1_combout ),
	.datad(!\Equal15~0_combout ),
	.datae(!\saved_read_data[9]~q ),
	.dataf(!\ctrl_wdata~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~16 .extended_lut = "off";
defparam \ctrl_wdata~16 .lut_mask = 64'h1111B1BB1F11BFBB;
defparam \ctrl_wdata~16 .shared_arith = "off";

dffeas \saved_read_data[10] (
	.clk(clk),
	.d(ctrl_rdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[10]~q ),
	.prn(vcc));
defparam \saved_read_data[10] .is_wysiwyg = "true";
defparam \saved_read_data[10] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~17 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~17 .extended_lut = "off";
defparam \ctrl_wdata~17 .lut_mask = 64'hFFFF7DF700000000;
defparam \ctrl_wdata~17 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~18 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_writedata_10),
	.datad(!\saved_read_data[10]~q ),
	.datae(!\ctrl_wdata~17_combout ),
	.dataf(!mif_rec_data_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~18 .extended_lut = "off";
defparam \ctrl_wdata~18 .lut_mask = 64'h03CF070703CF8F8F;
defparam \ctrl_wdata~18 .shared_arith = "off";

dffeas \saved_read_data[11] (
	.clk(clk),
	.d(ctrl_rdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[11]~q ),
	.prn(vcc));
defparam \saved_read_data[11] .is_wysiwyg = "true";
defparam \saved_read_data[11] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~19 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~19 .extended_lut = "off";
defparam \ctrl_wdata~19 .lut_mask = 64'hFFFF7FB700000000;
defparam \ctrl_wdata~19 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~20 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_writedata_11),
	.datad(!\saved_read_data[11]~q ),
	.datae(!\ctrl_wdata~19_combout ),
	.dataf(!mif_rec_data_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~20 .extended_lut = "off";
defparam \ctrl_wdata~20 .lut_mask = 64'h03CF070703CF8F8F;
defparam \ctrl_wdata~20 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~3 (
	.dataa(!uif_addr_offset_11),
	.datab(!\ctrl_next_state.CTRL_CHK_CHN~0_combout ),
	.datac(!\always6~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~3 .extended_lut = "off";
defparam \ctrl_addr~3 .lut_mask = 64'h3737373737373737;
defparam \ctrl_addr~3 .shared_arith = "off";

dffeas \saved_read_data[12] (
	.clk(clk),
	.d(ctrl_rdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[12]~q ),
	.prn(vcc));
defparam \saved_read_data[12] .is_wysiwyg = "true";
defparam \saved_read_data[12] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~21 (
	.dataa(!\mux_mif_addr[4]~0_combout ),
	.datab(!\mux_mif_addr[5]~1_combout ),
	.datac(!\mux_mif_addr[2]~2_combout ),
	.datad(!\mux_mif_addr[1]~3_combout ),
	.datae(!\Equal14~3_combout ),
	.dataf(!\Equal17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~21 .extended_lut = "off";
defparam \ctrl_wdata~21 .lut_mask = 64'hFFFF7F7700000000;
defparam \ctrl_wdata~21 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~22 (
	.dataa(!uif_ctrl_0),
	.datab(!uif_ctrl_1),
	.datac(!uif_writedata_12),
	.datad(!\saved_read_data[12]~q ),
	.datae(!\ctrl_wdata~21_combout ),
	.dataf(!mif_rec_data_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~22 .extended_lut = "off";
defparam \ctrl_wdata~22 .lut_mask = 64'h03CF070703CF8F8F;
defparam \ctrl_wdata~22 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~0 (
	.dataa(!\mux_mif_addr[1]~3_combout ),
	.datab(!\mux_mif_addr[0]~4_combout ),
	.datac(!\mux_mif_addr[3]~5_combout ),
	.datad(!\Equal14~0_combout ),
	.datae(!\Equal14~1_combout ),
	.dataf(!\Equal14~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'h0000000000000040;
defparam \Equal16~0 .shared_arith = "off";

dffeas \saved_read_data[13] (
	.clk(clk),
	.d(ctrl_rdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[13]~q ),
	.prn(vcc));
defparam \saved_read_data[13] .is_wysiwyg = "true";
defparam \saved_read_data[13] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~23 (
	.dataa(!uif_writedata_13),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!mif_rec_data_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~23 .extended_lut = "off";
defparam \ctrl_wdata~23 .lut_mask = 64'h4747474747474747;
defparam \ctrl_wdata~23 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~24 (
	.dataa(!uif_ctrl_1),
	.datab(!\Equal14~4_combout ),
	.datac(!\Equal16~0_combout ),
	.datad(!\Equal17~1_combout ),
	.datae(!\saved_read_data[13]~q ),
	.dataf(!\ctrl_wdata~23_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~24 .extended_lut = "off";
defparam \ctrl_wdata~24 .lut_mask = 64'h000002AAFD55FFFF;
defparam \ctrl_wdata~24 .shared_arith = "off";

dffeas \saved_read_data[14] (
	.clk(clk),
	.d(ctrl_rdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[14]~q ),
	.prn(vcc));
defparam \saved_read_data[14] .is_wysiwyg = "true";
defparam \saved_read_data[14] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~25 (
	.dataa(!uif_writedata_14),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!mif_rec_data_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~25 .extended_lut = "off";
defparam \ctrl_wdata~25 .lut_mask = 64'h4747474747474747;
defparam \ctrl_wdata~25 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~26 (
	.dataa(!uif_ctrl_1),
	.datab(!\Equal14~4_combout ),
	.datac(!\Equal16~0_combout ),
	.datad(!\Equal17~1_combout ),
	.datae(!\saved_read_data[14]~q ),
	.dataf(!\ctrl_wdata~25_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~26 .extended_lut = "off";
defparam \ctrl_wdata~26 .lut_mask = 64'h000002AAFD55FFFF;
defparam \ctrl_wdata~26 .shared_arith = "off";

dffeas \saved_read_data[15] (
	.clk(clk),
	.d(ctrl_rdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\saved_read_data[15]~q ),
	.prn(vcc));
defparam \saved_read_data[15] .is_wysiwyg = "true";
defparam \saved_read_data[15] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~27 (
	.dataa(!uif_writedata_15),
	.datab(!\ctrl_wdata~0_combout ),
	.datac(!mif_rec_data_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~27 .extended_lut = "off";
defparam \ctrl_wdata~27 .lut_mask = 64'h4747474747474747;
defparam \ctrl_wdata~27 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~28 (
	.dataa(!uif_ctrl_1),
	.datab(!\Equal14~4_combout ),
	.datac(!\Equal16~0_combout ),
	.datad(!\Equal17~1_combout ),
	.datae(!\saved_read_data[15]~q ),
	.dataf(!\ctrl_wdata~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~28 .extended_lut = "off";
defparam \ctrl_wdata~28 .lut_mask = 64'h000002AAFD55FFFF;
defparam \ctrl_wdata~28 .shared_arith = "off";

cyclonev_lcell_comb \mif_addr_mode~0 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_writedata_1),
	.datac(!uif_addr_offset_1),
	.datad(!uif_addr_offset_2),
	.datae(!\always0~0_combout ),
	.dataf(!mif_addr_mode1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_addr_mode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_addr_mode~0 .extended_lut = "off";
defparam \mif_addr_mode~0 .lut_mask = 64'h00001000FFFFBFFF;
defparam \mif_addr_mode~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_offset_cancellation (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	reconfig_mgmt_readdata_8,
	offset_cancellation_readdata_8,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write,
	grant_0,
	req_and_use_mutex,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	Equal0,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	offset_cancellation_done,
	ifsel_notdone_resync,
	comb,
	mutex_grant,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_write_data_1,
	master_write_data_2,
	master_write_data_0,
	master_write_data_3,
	master_write_data_4,
	master_write_data_5,
	master_write_data_6,
	master_write_data_7,
	master_write_data_8,
	master_write_data_9,
	master_write_data_10,
	master_write_data_11,
	master_write_data_12,
	master_write_data_13,
	master_write_data_14,
	master_write_data_15,
	out_narrow_0,
	out_narrow_1,
	out_narrow_2,
	out_narrow_3,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	reconfig_mgmt_readdata_8;
output 	offset_cancellation_readdata_8;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write;
input 	grant_0;
output 	req_and_use_mutex;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	Equal0;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
output 	offset_cancellation_done;
input 	ifsel_notdone_resync;
input 	comb;
output 	mutex_grant;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_write_data_1;
output 	master_write_data_2;
output 	master_write_data_0;
output 	master_write_data_3;
output 	master_write_data_4;
output 	master_write_data_5;
output 	master_write_data_6;
output 	master_write_data_7;
output 	master_write_data_8;
output 	master_write_data_9;
output 	master_write_data_10;
output 	master_write_data_11;
output 	master_write_data_12;
output 	master_write_data_13;
output 	master_write_data_14;
output 	master_write_data_15;
input 	out_narrow_0;
input 	out_narrow_1;
input 	out_narrow_2;
input 	out_narrow_3;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



RECONFIGURE_IP_alt_xcvr_reconfig_offset_cancellation_av offset_cancellation_av(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.reconfig_mgmt_readdata_8(reconfig_mgmt_readdata_8),
	.offset_cancellation_readdata_8(offset_cancellation_readdata_8),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.master_write1(master_write),
	.grant_0(grant_0),
	.req_and_use_mutex1(req_and_use_mutex),
	.master_address_2(master_address_2),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read1(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.Equal0(Equal0),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg(launch_reg),
	.wait_reg(wait_reg),
	.offset_cancellation_done(offset_cancellation_done),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.comb(comb),
	.mutex_grant(mutex_grant),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.master_write_data_1(master_write_data_1),
	.master_write_data_2(master_write_data_2),
	.master_write_data_0(master_write_data_0),
	.master_write_data_3(master_write_data_3),
	.master_write_data_4(master_write_data_4),
	.master_write_data_5(master_write_data_5),
	.master_write_data_6(master_write_data_6),
	.master_write_data_7(master_write_data_7),
	.master_write_data_8(master_write_data_8),
	.master_write_data_9(master_write_data_9),
	.master_write_data_10(master_write_data_10),
	.master_write_data_11(master_write_data_11),
	.master_write_data_12(master_write_data_12),
	.master_write_data_13(master_write_data_13),
	.master_write_data_14(master_write_data_14),
	.master_write_data_15(master_write_data_15),
	.out_narrow_0(out_narrow_0),
	.out_narrow_1(out_narrow_1),
	.out_narrow_2(out_narrow_2),
	.out_narrow_3(out_narrow_3),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0));

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_offset_cancellation_av (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	reconfig_mgmt_readdata_8,
	offset_cancellation_readdata_8,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write1,
	grant_0,
	req_and_use_mutex1,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read1,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	Equal0,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	offset_cancellation_done,
	ifsel_notdone_resync,
	comb,
	mutex_grant,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_write_data_1,
	master_write_data_2,
	master_write_data_0,
	master_write_data_3,
	master_write_data_4,
	master_write_data_5,
	master_write_data_6,
	master_write_data_7,
	master_write_data_8,
	master_write_data_9,
	master_write_data_10,
	master_write_data_11,
	master_write_data_12,
	master_write_data_13,
	master_write_data_14,
	master_write_data_15,
	out_narrow_0,
	out_narrow_1,
	out_narrow_2,
	out_narrow_3,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	reconfig_mgmt_readdata_8;
output 	offset_cancellation_readdata_8;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write1;
input 	grant_0;
output 	req_and_use_mutex1;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read1;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	Equal0;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
output 	offset_cancellation_done;
input 	ifsel_notdone_resync;
input 	comb;
output 	mutex_grant;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
input 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_write_data_1;
output 	master_write_data_2;
output 	master_write_data_0;
output 	master_write_data_3;
output 	master_write_data_4;
output 	master_write_data_5;
output 	master_write_data_6;
output 	master_write_data_7;
output 	master_write_data_8;
output 	master_write_data_9;
output 	master_write_data_10;
output 	master_write_data_11;
output 	master_write_data_12;
output 	master_write_data_13;
output 	master_write_data_14;
output 	master_write_data_15;
input 	out_narrow_0;
input 	out_narrow_1;
input 	out_narrow_2;
input 	out_narrow_3;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_cal_inst|alt_cal_busy~q ;
wire \alt_cal_inst|write_reg~q ;
wire \alt_cal_inst|read~q ;
wire \alt_cal_inst|alt_cal_channel[9]~q ;
wire \alt_cal_inst|alt_cal_channel[6]~q ;
wire \alt_cal_inst|alt_cal_channel[7]~q ;
wire \alt_cal_inst|alt_cal_channel[8]~q ;
wire \alt_cal_inst|alt_cal_channel[0]~q ;
wire \alt_cal_inst|alt_cal_channel[1]~q ;
wire \alt_cal_inst|alt_cal_channel[2]~q ;
wire \alt_cal_inst|alt_cal_channel[3]~q ;
wire \alt_cal_inst|alt_cal_channel[4]~q ;
wire \alt_cal_inst|alt_cal_channel[5]~q ;
wire \alt_cal_remap_addr[2]~q ;
wire \alt_cal_remap_addr[7]~q ;
wire \alt_cal_remap_addr[10]~q ;
wire \alt_cal_remap_addr[8]~q ;
wire \alt_cal_remap_addr[9]~q ;
wire \alt_cal_remap_addr[1]~q ;
wire \alt_cal_remap_addr[0]~q ;
wire \alt_cal_remap_addr[11]~q ;
wire \alt_cal_remap_addr[3]~q ;
wire \alt_cal_remap_addr[4]~q ;
wire \alt_cal_remap_addr[5]~q ;
wire \alt_cal_remap_addr[6]~q ;
wire \alt_cal_inst|address[1]~q ;
wire \alt_cal_inst|address[0]~q ;
wire \alt_cal_inst|address[4]~q ;
wire \start~q ;
wire \start0q~q ;
wire \alt_cal_dprio_busy~q ;
wire \alt_cal_inst|dataout[1]~q ;
wire \alt_cal_inst|dataout[2]~q ;
wire \alt_cal_inst|dataout[0]~q ;
wire \alt_cal_inst|dataout[3]~q ;
wire \alt_cal_inst|dataout[4]~q ;
wire \alt_cal_inst|dataout[5]~q ;
wire \alt_cal_inst|dataout[6]~q ;
wire \alt_cal_inst|dataout[7]~q ;
wire \alt_cal_inst|dataout[8]~q ;
wire \alt_cal_inst|dataout[9]~q ;
wire \alt_cal_inst|dataout[10]~q ;
wire \alt_cal_inst|dataout[11]~q ;
wire \alt_cal_inst|dataout[12]~q ;
wire \alt_cal_inst|dataout[13]~q ;
wire \alt_cal_inst|dataout[14]~q ;
wire \alt_cal_inst|dataout[15]~q ;
wire \start~0_combout ;
wire \start~1_combout ;
wire \Selector80~0_combout ;
wire \alt_cal_remap_addr[8]~0_combout ;
wire \alt_cal_dprio_datain[14]~q ;
wire \alt_cal_dprio_datain[1]~q ;
wire \alt_cal_dprio_datain[0]~q ;
wire \alt_cal_dprio_datain[3]~q ;
wire \alt_cal_dprio_datain[4]~q ;
wire \alt_cal_dprio_datain[5]~q ;
wire \alt_cal_dprio_datain[6]~q ;
wire \alt_cal_dprio_datain[7]~q ;
wire \alt_cal_dprio_datain[8]~q ;
wire \alt_cal_dprio_datain[9]~q ;
wire \alt_cal_dprio_datain[10]~q ;
wire \alt_cal_dprio_datain[11]~q ;
wire \alt_cal_dprio_datain[12]~q ;
wire \alt_cal_dprio_datain[13]~q ;
wire \alt_cal_dprio_datain[15]~q ;
wire \offset_cancellation_readdata[8]~0_combout ;
wire \master_write~0_combout ;
wire \always1~0_combout ;
wire \Selector16~0_combout ;
wire \state.GET_TESTBUS_DATA_STATE~q ;
wire \state.SET_OC_CALEN_ADDR_STATE~q ;
wire \state.SET_OC_CALEN_DATA_STATE~q ;
wire \state.START_OC_CALEN_STATE~q ;
wire \master_write_data[15]~6_combout ;
wire \pmutex_acquired~0_combout ;
wire \pmutex_acquired~q ;
wire \Selector24~0_combout ;
wire \state.ADDRESS_OFFSET_STATE~q ;
wire \Selector14~0_combout ;
wire \write_read_control~0_combout ;
wire \write_read_control~q ;
wire \Selector17~0_combout ;
wire \state.WRITE_DATA_STATE~q ;
wire \Selector18~0_combout ;
wire \state.CONTROL_STATE~q ;
wire \state.BUSY_STATE~q ;
wire \state~46_combout ;
wire \state.WRITE_DONE_STATE~q ;
wire \Selector25~0_combout ;
wire \state.READ_DATA_STATE~q ;
wire \Selector29~0_combout ;
wire \Selector29~1_combout ;
wire \state.WAIT_FOR_NEXT_STATE~q ;
wire \Selector0~3_combout ;
wire \prev_logical_channel[9]~q ;
wire \Equal2~0_combout ;
wire \prev_logical_channel[6]~q ;
wire \prev_logical_channel[7]~q ;
wire \prev_logical_channel[8]~q ;
wire \Equal2~1_combout ;
wire \prev_logical_channel[0]~q ;
wire \prev_logical_channel[1]~q ;
wire \prev_logical_channel[2]~q ;
wire \Equal2~2_combout ;
wire \prev_logical_channel[3]~q ;
wire \prev_logical_channel[4]~q ;
wire \prev_logical_channel[5]~q ;
wire \Equal2~3_combout ;
wire \Selector45~7_combout ;
wire \Selector28~0_combout ;
wire \state.RELEASE_PMUTEX_STATE~q ;
wire \state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE~q ;
wire \state.RELEASE_PHY_RESET_OVERRIDE_DATA_STATE~q ;
wire \state.RELEASE_PHY_RESET_OVERRIDE_START_STATE~q ;
wire \state.RELEASE_OC_CALEN_DATA_STATE~q ;
wire \state.RELEASE_OC_CALEN_START_STATE~q ;
wire \state.RELEASE_OC_CALEN_DONE_STATE~q ;
wire \Selector15~0_combout ;
wire \Selector15~1_combout ;
wire \state.000000~q ;
wire \Selector16~1_combout ;
wire \Selector16~2_combout ;
wire \state.LOGICAL_ADDRESS_STATE~q ;
wire \state.READ_PHY_ADDR_STATE~q ;
wire \state~44_combout ;
wire \state.CHECK_PHY_ADDR_STATE~q ;
wire \Selector21~0_combout ;
wire \Selector21~1_combout ;
wire \state.SET_ADDR_OFFSET_REQ_STATE~q ;
wire \state.REQUEST_CONTROL_STATE~q ;
wire \Selector23~0_combout ;
wire \state.READ_REQ_DATA_STATE~q ;
wire \state~45_combout ;
wire \state.CHECK_REQ_DATA_STATE~q ;
wire \Selector26~0_combout ;
wire \state.ACQUIRE_PMUTEX_STATE~q ;
wire \Selector27~0_combout ;
wire \state.READ_PMUTEX_STATE~q ;
wire \state~43_combout ;
wire \state.CHECK_PMUTEX_STATE~q ;
wire \Selector38~0_combout ;
wire \Selector38~1_combout ;
wire \state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ;
wire \state.SET_PHY_RESET_OVERRIDE_DATA_STATE~q ;
wire \state.SET_PHY_RESET_OVERRIDE_START_STATE~q ;
wire \state.GET_TESTBUS_ADDR_STATE~q ;
wire \Selector78~0_combout ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \Selector1~3_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector0~2_combout ;
wire \Selector0~4_combout ;
wire \Selector0~5_combout ;
wire \Selector0~6_combout ;
wire \Selector0~7_combout ;
wire \offset_cancellation_done~2_combout ;
wire \master_address~0_combout ;
wire \Selector45~0_combout ;
wire \Selector44~0_combout ;
wire \WideOr2~0_combout ;
wire \Selector44~1_combout ;
wire \Selector44~2_combout ;
wire \Selector45~1_combout ;
wire \Selector45~2_combout ;
wire \Selector45~3_combout ;
wire \Selector44~4_combout ;
wire \Selector44~3_combout ;
wire \Selector46~0_combout ;
wire \Selector45~4_combout ;
wire \Selector46~1_combout ;
wire \Selector46~2_combout ;
wire \Selector46~3_combout ;
wire \Selector46~4_combout ;
wire \Selector46~5_combout ;
wire \Selector1~4_combout ;
wire \Selector46~6_combout ;
wire \Selector45~5_combout ;
wire \Selector45~6_combout ;
wire \Selector45~8_combout ;
wire \Selector45~9_combout ;
wire \Selector45~10_combout ;
wire \Selector45~11_combout ;
wire \Selector1~5_combout ;
wire \Selector1~6_combout ;
wire \WideOr34~0_combout ;
wire \Selector1~7_combout ;
wire \Selector1~8_combout ;
wire \Selector1~9_combout ;
wire \Selector1~10_combout ;
wire \oc_started~0_combout ;
wire \oc_started~q ;
wire \WideOr34~combout ;
wire \Selector67~0_combout ;
wire \Selector77~0_combout ;
wire \Selector77~1_combout ;
wire \Selector77~2_combout ;
wire \Selector77~3_combout ;
wire \Selector77~4_combout ;
wire \Selector77~5_combout ;
wire \Selector76~0_combout ;
wire \Selector76~1_combout ;
wire \Selector76~2_combout ;
wire \master_write_data[7]~0_combout ;
wire \Selector76~3_combout ;
wire \Selector76~4_combout ;
wire \Selector76~5_combout ;
wire \Selector78~1_combout ;
wire \Selector78~2_combout ;
wire \Selector78~3_combout ;
wire \Selector78~4_combout ;
wire \master_write_data[7]~1_combout ;
wire \Selector78~5_combout ;
wire \Selector78~6_combout ;
wire \Selector78~7_combout ;
wire \Selector75~0_combout ;
wire \Selector75~1_combout ;
wire \Selector75~2_combout ;
wire \Selector75~3_combout ;
wire \Selector75~4_combout ;
wire \Selector74~0_combout ;
wire \Selector74~1_combout ;
wire \Selector74~2_combout ;
wire \master_write_data[7]~2_combout ;
wire \Equal2~4_combout ;
wire \Selector73~0_combout ;
wire \master_write_data[7]~3_combout ;
wire \master_write_data[7]~4_combout ;
wire \Selector72~0_combout ;
wire \Selector71~0_combout ;
wire \Selector70~0_combout ;
wire \Selector69~0_combout ;
wire \Selector68~0_combout ;
wire \master_write_data[15]~5_combout ;
wire \master_write_data[15]~7_combout ;
wire \master_write_data[15]~8_combout ;
wire \master_write_data[15]~9_combout ;
wire \master_write_data[15]~10_combout ;
wire \Selector67~2_combout ;
wire \Selector67~1_combout ;
wire \Selector67~3_combout ;
wire \Selector66~0_combout ;
wire \master_write_data[12]~11_combout ;
wire \master_write_data[12]~12_combout ;
wire \master_write_data[12]~13_combout ;
wire \Selector65~0_combout ;
wire \Selector64~0_combout ;
wire \Selector63~0_combout ;


RECONFIGURE_IP_alt_arbiter_acq_3 mutex_inst(
	.grant_0(grant_0),
	.req_and_use_mutex(req_and_use_mutex1),
	.mutex_grant(mutex_grant));

RECONFIGURE_IP_alt_cal_av_1 alt_cal_inst(
	.alt_cal_busy1(\alt_cal_inst|alt_cal_busy~q ),
	.write_reg1(\alt_cal_inst|write_reg~q ),
	.read1(\alt_cal_inst|read~q ),
	.alt_cal_channel_9(\alt_cal_inst|alt_cal_channel[9]~q ),
	.alt_cal_channel_6(\alt_cal_inst|alt_cal_channel[6]~q ),
	.alt_cal_channel_7(\alt_cal_inst|alt_cal_channel[7]~q ),
	.alt_cal_channel_8(\alt_cal_inst|alt_cal_channel[8]~q ),
	.alt_cal_channel_0(\alt_cal_inst|alt_cal_channel[0]~q ),
	.alt_cal_channel_1(\alt_cal_inst|alt_cal_channel[1]~q ),
	.alt_cal_channel_2(\alt_cal_inst|alt_cal_channel[2]~q ),
	.alt_cal_channel_3(\alt_cal_inst|alt_cal_channel[3]~q ),
	.alt_cal_channel_4(\alt_cal_inst|alt_cal_channel[4]~q ),
	.alt_cal_channel_5(\alt_cal_inst|alt_cal_channel[5]~q ),
	.alt_cal_remap_addr_2(\alt_cal_remap_addr[2]~q ),
	.alt_cal_remap_addr_7(\alt_cal_remap_addr[7]~q ),
	.alt_cal_remap_addr_10(\alt_cal_remap_addr[10]~q ),
	.alt_cal_remap_addr_8(\alt_cal_remap_addr[8]~q ),
	.alt_cal_remap_addr_9(\alt_cal_remap_addr[9]~q ),
	.alt_cal_remap_addr_1(\alt_cal_remap_addr[1]~q ),
	.alt_cal_remap_addr_0(\alt_cal_remap_addr[0]~q ),
	.alt_cal_remap_addr_11(\alt_cal_remap_addr[11]~q ),
	.alt_cal_remap_addr_3(\alt_cal_remap_addr[3]~q ),
	.alt_cal_remap_addr_4(\alt_cal_remap_addr[4]~q ),
	.alt_cal_remap_addr_5(\alt_cal_remap_addr[5]~q ),
	.alt_cal_remap_addr_6(\alt_cal_remap_addr[6]~q ),
	.address_1(\alt_cal_inst|address[1]~q ),
	.address_0(\alt_cal_inst|address[0]~q ),
	.address_4(\alt_cal_inst|address[4]~q ),
	.reset(ifsel_notdone_resync),
	.start(\start~q ),
	.start0q(\start0q~q ),
	.alt_cal_dprio_busy(\alt_cal_dprio_busy~q ),
	.dataout_1(\alt_cal_inst|dataout[1]~q ),
	.dataout_2(\alt_cal_inst|dataout[2]~q ),
	.dataout_0(\alt_cal_inst|dataout[0]~q ),
	.dataout_3(\alt_cal_inst|dataout[3]~q ),
	.dataout_4(\alt_cal_inst|dataout[4]~q ),
	.dataout_5(\alt_cal_inst|dataout[5]~q ),
	.dataout_6(\alt_cal_inst|dataout[6]~q ),
	.dataout_7(\alt_cal_inst|dataout[7]~q ),
	.dataout_8(\alt_cal_inst|dataout[8]~q ),
	.dataout_9(\alt_cal_inst|dataout[9]~q ),
	.dataout_10(\alt_cal_inst|dataout[10]~q ),
	.dataout_11(\alt_cal_inst|dataout[11]~q ),
	.dataout_12(\alt_cal_inst|dataout[12]~q ),
	.dataout_13(\alt_cal_inst|dataout[13]~q ),
	.dataout_14(\alt_cal_inst|dataout[14]~q ),
	.dataout_15(\alt_cal_inst|dataout[15]~q ),
	.alt_cal_dprio_datain_14(\alt_cal_dprio_datain[14]~q ),
	.alt_cal_dprio_datain_1(\alt_cal_dprio_datain[1]~q ),
	.alt_cal_dprio_datain_0(\alt_cal_dprio_datain[0]~q ),
	.alt_cal_dprio_datain_3(\alt_cal_dprio_datain[3]~q ),
	.alt_cal_dprio_datain_4(\alt_cal_dprio_datain[4]~q ),
	.alt_cal_dprio_datain_5(\alt_cal_dprio_datain[5]~q ),
	.alt_cal_dprio_datain_6(\alt_cal_dprio_datain[6]~q ),
	.alt_cal_dprio_datain_7(\alt_cal_dprio_datain[7]~q ),
	.alt_cal_dprio_datain_8(\alt_cal_dprio_datain[8]~q ),
	.alt_cal_dprio_datain_9(\alt_cal_dprio_datain[9]~q ),
	.alt_cal_dprio_datain_10(\alt_cal_dprio_datain[10]~q ),
	.alt_cal_dprio_datain_11(\alt_cal_dprio_datain[11]~q ),
	.alt_cal_dprio_datain_12(\alt_cal_dprio_datain[12]~q ),
	.alt_cal_dprio_datain_13(\alt_cal_dprio_datain[13]~q ),
	.alt_cal_dprio_datain_15(\alt_cal_dprio_datain[15]~q ),
	.out_narrow_0(out_narrow_0),
	.out_narrow_1(out_narrow_1),
	.out_narrow_2(out_narrow_2),
	.out_narrow_3(out_narrow_3),
	.clock(mgmt_clk_clk));

RECONFIGURE_IP_altera_wait_generate_2 wait_gen(
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg1(launch_reg),
	.wait_reg1(wait_reg),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.launch_signal(comb),
	.mgmt_clk_clk(mgmt_clk_clk));

dffeas \alt_cal_remap_addr[2] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_2),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[2]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[2] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[2] .power_up = "low";

dffeas \alt_cal_remap_addr[7] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_7),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[7]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[7] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[7] .power_up = "low";

dffeas \alt_cal_remap_addr[10] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_10),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[10]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[10] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[10] .power_up = "low";

dffeas \alt_cal_remap_addr[8] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_8),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[8]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[8] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[8] .power_up = "low";

dffeas \alt_cal_remap_addr[9] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_9),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[9]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[9] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[9] .power_up = "low";

dffeas \alt_cal_remap_addr[1] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_1),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[1]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[1] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[1] .power_up = "low";

dffeas \alt_cal_remap_addr[0] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_0),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[0]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[0] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[0] .power_up = "low";

dffeas \alt_cal_remap_addr[11] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_11),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[11]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[11] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[11] .power_up = "low";

dffeas \alt_cal_remap_addr[3] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_3),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[3]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[3] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[3] .power_up = "low";

dffeas \alt_cal_remap_addr[4] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_4),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[4]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[4] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[4] .power_up = "low";

dffeas \alt_cal_remap_addr[5] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_5),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[5]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[5] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[5] .power_up = "low";

dffeas \alt_cal_remap_addr[6] (
	.clk(mgmt_clk_clk),
	.d(\WideOr2~0_combout ),
	.asdata(basic_reconfig_readdata_6),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Selector21~0_combout ),
	.ena(\alt_cal_remap_addr[8]~0_combout ),
	.q(\alt_cal_remap_addr[6]~q ),
	.prn(vcc));
defparam \alt_cal_remap_addr[6] .is_wysiwyg = "true";
defparam \alt_cal_remap_addr[6] .power_up = "low";

dffeas start(
	.clk(mgmt_clk_clk),
	.d(\start~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start~1_combout ),
	.q(\start~q ),
	.prn(vcc));
defparam start.is_wysiwyg = "true";
defparam start.power_up = "low";

dffeas start0q(
	.clk(mgmt_clk_clk),
	.d(\start~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start~1_combout ),
	.q(\start0q~q ),
	.prn(vcc));
defparam start0q.is_wysiwyg = "true";
defparam start0q.power_up = "low";

dffeas alt_cal_dprio_busy(
	.clk(mgmt_clk_clk),
	.d(\Selector80~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\alt_cal_dprio_busy~q ),
	.prn(vcc));
defparam alt_cal_dprio_busy.is_wysiwyg = "true";
defparam alt_cal_dprio_busy.power_up = "low";

cyclonev_lcell_comb \start~0 (
	.dataa(!Equal0),
	.datab(!reconfig_mgmt_readdata_8),
	.datac(!reconfig_mgmt_write),
	.datad(!reconfig_mgmt_writedata_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\start~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \start~0 .extended_lut = "off";
defparam \start~0 .lut_mask = 64'h0001000100010001;
defparam \start~0 .shared_arith = "off";

cyclonev_lcell_comb \start~1 (
	.dataa(!Equal0),
	.datab(!reconfig_mgmt_readdata_8),
	.datac(!reconfig_mgmt_read),
	.datad(!reconfig_mgmt_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\start~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \start~1 .extended_lut = "off";
defparam \start~1 .lut_mask = 64'hFABAFABAFABAFABA;
defparam \start~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector80~0 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.READ_DATA_STATE~q ),
	.datac(!\state.BUSY_STATE~q ),
	.datad(!\alt_cal_dprio_busy~q ),
	.datae(!\state.WRITE_DONE_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector80~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector80~0 .extended_lut = "off";
defparam \Selector80~0 .lut_mask = 64'h0FEF0F2F0FEF0F2F;
defparam \Selector80~0 .shared_arith = "off";

cyclonev_lcell_comb \alt_cal_remap_addr[8]~0 (
	.dataa(!basic_reconfig_readdata_2),
	.datab(!\state.000000~q ),
	.datac(!\state.CHECK_PHY_ADDR_STATE~q ),
	.datad(!\state.CHECK_REQ_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\alt_cal_remap_addr[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \alt_cal_remap_addr[8]~0 .extended_lut = "off";
defparam \alt_cal_remap_addr[8]~0 .lut_mask = 64'hCFAACFAACFAACFAA;
defparam \alt_cal_remap_addr[8]~0 .shared_arith = "off";

dffeas \alt_cal_dprio_datain[14] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_14),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[14]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[14] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[14] .power_up = "low";

dffeas \alt_cal_dprio_datain[1] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[1]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[1] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[1] .power_up = "low";

dffeas \alt_cal_dprio_datain[0] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[0]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[0] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[0] .power_up = "low";

dffeas \alt_cal_dprio_datain[3] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[3]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[3] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[3] .power_up = "low";

dffeas \alt_cal_dprio_datain[4] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[4]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[4] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[4] .power_up = "low";

dffeas \alt_cal_dprio_datain[5] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[5]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[5] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[5] .power_up = "low";

dffeas \alt_cal_dprio_datain[6] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[6]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[6] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[6] .power_up = "low";

dffeas \alt_cal_dprio_datain[7] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[7]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[7] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[7] .power_up = "low";

dffeas \alt_cal_dprio_datain[8] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[8]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[8] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[8] .power_up = "low";

dffeas \alt_cal_dprio_datain[9] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[9]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[9] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[9] .power_up = "low";

dffeas \alt_cal_dprio_datain[10] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_10),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[10]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[10] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[10] .power_up = "low";

dffeas \alt_cal_dprio_datain[11] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_11),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[11]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[11] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[11] .power_up = "low";

dffeas \alt_cal_dprio_datain[12] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_12),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[12]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[12] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[12] .power_up = "low";

dffeas \alt_cal_dprio_datain[13] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_13),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[13]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[13] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[13] .power_up = "low";

dffeas \alt_cal_dprio_datain[15] (
	.clk(mgmt_clk_clk),
	.d(basic_reconfig_readdata_15),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector29~0_combout ),
	.q(\alt_cal_dprio_datain[15]~q ),
	.prn(vcc));
defparam \alt_cal_dprio_datain[15] .is_wysiwyg = "true";
defparam \alt_cal_dprio_datain[15] .power_up = "low";

dffeas \offset_cancellation_readdata[8] (
	.clk(mgmt_clk_clk),
	.d(\offset_cancellation_readdata[8]~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(offset_cancellation_readdata_8),
	.prn(vcc));
defparam \offset_cancellation_readdata[8] .is_wysiwyg = "true";
defparam \offset_cancellation_readdata[8] .power_up = "low";

dffeas master_write(
	.clk(mgmt_clk_clk),
	.d(\Selector0~7_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write1),
	.prn(vcc));
defparam master_write.is_wysiwyg = "true";
defparam master_write.power_up = "low";

dffeas req_and_use_mutex(
	.clk(mgmt_clk_clk),
	.d(\offset_cancellation_done~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(req_and_use_mutex1),
	.prn(vcc));
defparam req_and_use_mutex.is_wysiwyg = "true";
defparam req_and_use_mutex.power_up = "low";

dffeas \master_address[2] (
	.clk(mgmt_clk_clk),
	.d(\Selector44~3_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_2),
	.prn(vcc));
defparam \master_address[2] .is_wysiwyg = "true";
defparam \master_address[2] .power_up = "low";

dffeas \master_address[0] (
	.clk(mgmt_clk_clk),
	.d(\Selector46~6_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_0),
	.prn(vcc));
defparam \master_address[0] .is_wysiwyg = "true";
defparam \master_address[0] .power_up = "low";

dffeas \master_address[1] (
	.clk(mgmt_clk_clk),
	.d(\Selector45~11_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_1),
	.prn(vcc));
defparam \master_address[1] .is_wysiwyg = "true";
defparam \master_address[1] .power_up = "low";

dffeas master_read(
	.clk(mgmt_clk_clk),
	.d(\Selector1~10_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_read1),
	.prn(vcc));
defparam master_read.is_wysiwyg = "true";
defparam master_read.power_up = "low";

cyclonev_lcell_comb \offset_cancellation_done~1 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.000000~q ),
	.datac(!\oc_started~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(offset_cancellation_done),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_cancellation_done~1 .extended_lut = "off";
defparam \offset_cancellation_done~1 .lut_mask = 64'h0808080808080808;
defparam \offset_cancellation_done~1 .shared_arith = "off";

dffeas \master_write_data[1] (
	.clk(mgmt_clk_clk),
	.d(\Selector77~5_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write_data_1),
	.prn(vcc));
defparam \master_write_data[1] .is_wysiwyg = "true";
defparam \master_write_data[1] .power_up = "low";

dffeas \master_write_data[2] (
	.clk(mgmt_clk_clk),
	.d(\Selector76~5_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write_data_2),
	.prn(vcc));
defparam \master_write_data[2] .is_wysiwyg = "true";
defparam \master_write_data[2] .power_up = "low";

dffeas \master_write_data[0] (
	.clk(mgmt_clk_clk),
	.d(\Selector78~7_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write_data_0),
	.prn(vcc));
defparam \master_write_data[0] .is_wysiwyg = "true";
defparam \master_write_data[0] .power_up = "low";

dffeas \master_write_data[3] (
	.clk(mgmt_clk_clk),
	.d(\Selector75~4_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write_data_3),
	.prn(vcc));
defparam \master_write_data[3] .is_wysiwyg = "true";
defparam \master_write_data[3] .power_up = "low";

dffeas \master_write_data[4] (
	.clk(mgmt_clk_clk),
	.d(\Selector74~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write_data_4),
	.prn(vcc));
defparam \master_write_data[4] .is_wysiwyg = "true";
defparam \master_write_data[4] .power_up = "low";

dffeas \master_write_data[5] (
	.clk(mgmt_clk_clk),
	.d(\Selector73~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[7]~4_combout ),
	.q(master_write_data_5),
	.prn(vcc));
defparam \master_write_data[5] .is_wysiwyg = "true";
defparam \master_write_data[5] .power_up = "low";

dffeas \master_write_data[6] (
	.clk(mgmt_clk_clk),
	.d(\Selector72~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[7]~4_combout ),
	.q(master_write_data_6),
	.prn(vcc));
defparam \master_write_data[6] .is_wysiwyg = "true";
defparam \master_write_data[6] .power_up = "low";

dffeas \master_write_data[7] (
	.clk(mgmt_clk_clk),
	.d(\Selector71~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[7]~4_combout ),
	.q(master_write_data_7),
	.prn(vcc));
defparam \master_write_data[7] .is_wysiwyg = "true";
defparam \master_write_data[7] .power_up = "low";

dffeas \master_write_data[8] (
	.clk(mgmt_clk_clk),
	.d(\Selector70~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[7]~4_combout ),
	.q(master_write_data_8),
	.prn(vcc));
defparam \master_write_data[8] .is_wysiwyg = "true";
defparam \master_write_data[8] .power_up = "low";

dffeas \master_write_data[9] (
	.clk(mgmt_clk_clk),
	.d(\Selector69~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[7]~4_combout ),
	.q(master_write_data_9),
	.prn(vcc));
defparam \master_write_data[9] .is_wysiwyg = "true";
defparam \master_write_data[9] .power_up = "low";

dffeas \master_write_data[10] (
	.clk(mgmt_clk_clk),
	.d(\Selector68~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[15]~10_combout ),
	.q(master_write_data_10),
	.prn(vcc));
defparam \master_write_data[10] .is_wysiwyg = "true";
defparam \master_write_data[10] .power_up = "low";

dffeas \master_write_data[11] (
	.clk(mgmt_clk_clk),
	.d(\Selector67~3_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write_data_11),
	.prn(vcc));
defparam \master_write_data[11] .is_wysiwyg = "true";
defparam \master_write_data[11] .power_up = "low";

dffeas \master_write_data[12] (
	.clk(mgmt_clk_clk),
	.d(\Selector66~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[12]~13_combout ),
	.q(master_write_data_12),
	.prn(vcc));
defparam \master_write_data[12] .is_wysiwyg = "true";
defparam \master_write_data[12] .power_up = "low";

dffeas \master_write_data[13] (
	.clk(mgmt_clk_clk),
	.d(\Selector65~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[12]~13_combout ),
	.q(master_write_data_13),
	.prn(vcc));
defparam \master_write_data[13] .is_wysiwyg = "true";
defparam \master_write_data[13] .power_up = "low";

dffeas \master_write_data[14] (
	.clk(mgmt_clk_clk),
	.d(\Selector64~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[15]~10_combout ),
	.q(master_write_data_14),
	.prn(vcc));
defparam \master_write_data[14] .is_wysiwyg = "true";
defparam \master_write_data[14] .power_up = "low";

dffeas \master_write_data[15] (
	.clk(mgmt_clk_clk),
	.d(\Selector63~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write_data[15]~10_combout ),
	.q(master_write_data_15),
	.prn(vcc));
defparam \master_write_data[15] .is_wysiwyg = "true";
defparam \master_write_data[15] .power_up = "low";

cyclonev_lcell_comb \offset_cancellation_readdata[8]~0 (
	.dataa(!offset_cancellation_readdata_8),
	.datab(!reconfig_mgmt_readdata_8),
	.datac(!comb),
	.datad(!\alt_cal_inst|alt_cal_busy~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_cancellation_readdata[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_cancellation_readdata[8]~0 .extended_lut = "off";
defparam \offset_cancellation_readdata[8]~0 .lut_mask = 64'h5457545754575457;
defparam \offset_cancellation_readdata[8]~0 .shared_arith = "off";

cyclonev_lcell_comb \master_write~0 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write~0 .extended_lut = "off";
defparam \master_write~0 .lut_mask = 64'h0404040404040404;
defparam \master_write~0 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!\alt_cal_inst|write_reg~q ),
	.datab(!\alt_cal_inst|read~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'h8888888888888888;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'h1111111111111111;
defparam \Selector16~0 .shared_arith = "off";

dffeas \state.GET_TESTBUS_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.GET_TESTBUS_ADDR_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.GET_TESTBUS_DATA_STATE~q ),
	.prn(vcc));
defparam \state.GET_TESTBUS_DATA_STATE .is_wysiwyg = "true";
defparam \state.GET_TESTBUS_DATA_STATE .power_up = "low";

dffeas \state.SET_OC_CALEN_ADDR_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.GET_TESTBUS_DATA_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.SET_OC_CALEN_ADDR_STATE~q ),
	.prn(vcc));
defparam \state.SET_OC_CALEN_ADDR_STATE .is_wysiwyg = "true";
defparam \state.SET_OC_CALEN_ADDR_STATE .power_up = "low";

dffeas \state.SET_OC_CALEN_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.SET_OC_CALEN_ADDR_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.SET_OC_CALEN_DATA_STATE~q ),
	.prn(vcc));
defparam \state.SET_OC_CALEN_DATA_STATE .is_wysiwyg = "true";
defparam \state.SET_OC_CALEN_DATA_STATE .power_up = "low";

dffeas \state.START_OC_CALEN_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.SET_OC_CALEN_DATA_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.START_OC_CALEN_STATE~q ),
	.prn(vcc));
defparam \state.START_OC_CALEN_STATE .is_wysiwyg = "true";
defparam \state.START_OC_CALEN_STATE .power_up = "low";

cyclonev_lcell_comb \master_write_data[15]~6 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest1),
	.datac(!lif_waitrequest),
	.datad(!basic_reconfig_waitrequest),
	.datae(!lif_waitrequest2),
	.dataf(!\state.RELEASE_PMUTEX_STATE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[15]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[15]~6 .extended_lut = "off";
defparam \master_write_data[15]~6 .lut_mask = 64'h0000000040000000;
defparam \master_write_data[15]~6 .shared_arith = "off";

cyclonev_lcell_comb \pmutex_acquired~0 (
	.dataa(!\state.RELEASE_PMUTEX_STATE~q ),
	.datab(!\Selector38~0_combout ),
	.datac(!\pmutex_acquired~q ),
	.datad(!\master_write_data[15]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pmutex_acquired~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pmutex_acquired~0 .extended_lut = "off";
defparam \pmutex_acquired~0 .lut_mask = 64'h2F222F222F222F22;
defparam \pmutex_acquired~0 .shared_arith = "off";

dffeas pmutex_acquired(
	.clk(mgmt_clk_clk),
	.d(\pmutex_acquired~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pmutex_acquired~q ),
	.prn(vcc));
defparam pmutex_acquired.is_wysiwyg = "true";
defparam pmutex_acquired.power_up = "low";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!basic_reconfig_readdata_2),
	.datab(!\master_write~0_combout ),
	.datac(!\state.START_OC_CALEN_STATE~q ),
	.datad(!\state.ADDRESS_OFFSET_STATE~q ),
	.datae(!\state.CHECK_REQ_DATA_STATE~q ),
	.dataf(!\pmutex_acquired~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h03CF03CF03CF57DF;
defparam \Selector24~0 .shared_arith = "off";

dffeas \state.ADDRESS_OFFSET_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ADDRESS_OFFSET_STATE~q ),
	.prn(vcc));
defparam \state.ADDRESS_OFFSET_STATE .is_wysiwyg = "true";
defparam \state.ADDRESS_OFFSET_STATE .power_up = "low";

cyclonev_lcell_comb \Selector14~0 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.000000~q ),
	.datac(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~0 .extended_lut = "off";
defparam \Selector14~0 .lut_mask = 64'h3232323232323232;
defparam \Selector14~0 .shared_arith = "off";

cyclonev_lcell_comb \write_read_control~0 (
	.dataa(!\alt_cal_inst|write_reg~q ),
	.datab(!\alt_cal_inst|read~q ),
	.datac(!\write_read_control~q ),
	.datad(!\Selector14~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_read_control~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_read_control~0 .extended_lut = "off";
defparam \write_read_control~0 .lut_mask = 64'h5D0F5D0F5D0F5D0F;
defparam \write_read_control~0 .shared_arith = "off";

dffeas write_read_control(
	.clk(mgmt_clk_clk),
	.d(\write_read_control~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write_read_control~q ),
	.prn(vcc));
defparam write_read_control.is_wysiwyg = "true";
defparam write_read_control.power_up = "low";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!\state.ADDRESS_OFFSET_STATE~q ),
	.datab(!\write_read_control~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'h1111111111111111;
defparam \Selector17~0 .shared_arith = "off";

dffeas \state.WRITE_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.WRITE_DATA_STATE~q ),
	.prn(vcc));
defparam \state.WRITE_DATA_STATE .is_wysiwyg = "true";
defparam \state.WRITE_DATA_STATE .power_up = "low";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.CONTROL_STATE~q ),
	.datac(!\state.WRITE_DATA_STATE~q ),
	.datad(!\state.ADDRESS_OFFSET_STATE~q ),
	.datae(!\write_read_control~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h2777272727772727;
defparam \Selector18~0 .shared_arith = "off";

dffeas \state.CONTROL_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CONTROL_STATE~q ),
	.prn(vcc));
defparam \state.CONTROL_STATE .is_wysiwyg = "true";
defparam \state.CONTROL_STATE .power_up = "low";

dffeas \state.BUSY_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.CONTROL_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.BUSY_STATE~q ),
	.prn(vcc));
defparam \state.BUSY_STATE .is_wysiwyg = "true";
defparam \state.BUSY_STATE .power_up = "low";

cyclonev_lcell_comb \state~46 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.BUSY_STATE~q ),
	.datac(!\write_read_control~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~46 .extended_lut = "off";
defparam \state~46 .lut_mask = 64'h0101010101010101;
defparam \state~46 .shared_arith = "off";

dffeas \state.WRITE_DONE_STATE (
	.clk(mgmt_clk_clk),
	.d(\state~46_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.WRITE_DONE_STATE~q ),
	.prn(vcc));
defparam \state.WRITE_DONE_STATE .is_wysiwyg = "true";
defparam \state.WRITE_DONE_STATE .power_up = "low";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!\state.BUSY_STATE~q ),
	.datab(!\write_read_control~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h4444444444444444;
defparam \Selector25~0 .shared_arith = "off";

dffeas \state.READ_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.READ_DATA_STATE~q ),
	.prn(vcc));
defparam \state.READ_DATA_STATE .is_wysiwyg = "true";
defparam \state.READ_DATA_STATE .power_up = "low";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest1),
	.datac(!lif_waitrequest),
	.datad(!basic_reconfig_waitrequest),
	.datae(!lif_waitrequest2),
	.dataf(!\state.READ_DATA_STATE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'h0000000040000000;
defparam \Selector29~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~1 (
	.dataa(!\always1~0_combout ),
	.datab(!\Selector16~0_combout ),
	.datac(!\state.WRITE_DONE_STATE~q ),
	.datad(!\Selector29~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~1 .extended_lut = "off";
defparam \Selector29~1 .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \Selector29~1 .shared_arith = "off";

dffeas \state.WAIT_FOR_NEXT_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector29~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.WAIT_FOR_NEXT_STATE~q ),
	.prn(vcc));
defparam \state.WAIT_FOR_NEXT_STATE .is_wysiwyg = "true";
defparam \state.WAIT_FOR_NEXT_STATE .power_up = "low";

cyclonev_lcell_comb \Selector0~3 (
	.dataa(!\state.000000~q ),
	.datab(!\alt_cal_inst|write_reg~q ),
	.datac(!\alt_cal_inst|read~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~3 .extended_lut = "off";
defparam \Selector0~3 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \Selector0~3 .shared_arith = "off";

dffeas \prev_logical_channel[9] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[9]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[9]~q ),
	.prn(vcc));
defparam \prev_logical_channel[9] .is_wysiwyg = "true";
defparam \prev_logical_channel[9] .power_up = "low";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!\prev_logical_channel[9]~q ),
	.datab(!\alt_cal_inst|alt_cal_channel[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h6666666666666666;
defparam \Equal2~0 .shared_arith = "off";

dffeas \prev_logical_channel[6] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[6]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[6]~q ),
	.prn(vcc));
defparam \prev_logical_channel[6] .is_wysiwyg = "true";
defparam \prev_logical_channel[6] .power_up = "low";

dffeas \prev_logical_channel[7] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[7]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[7]~q ),
	.prn(vcc));
defparam \prev_logical_channel[7] .is_wysiwyg = "true";
defparam \prev_logical_channel[7] .power_up = "low";

dffeas \prev_logical_channel[8] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[8]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[8]~q ),
	.prn(vcc));
defparam \prev_logical_channel[8] .is_wysiwyg = "true";
defparam \prev_logical_channel[8] .power_up = "low";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!\prev_logical_channel[6]~q ),
	.datab(!\alt_cal_inst|alt_cal_channel[6]~q ),
	.datac(!\prev_logical_channel[7]~q ),
	.datad(!\alt_cal_inst|alt_cal_channel[7]~q ),
	.datae(!\prev_logical_channel[8]~q ),
	.dataf(!\alt_cal_inst|alt_cal_channel[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'h9009000000009009;
defparam \Equal2~1 .shared_arith = "off";

dffeas \prev_logical_channel[0] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[0]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[0]~q ),
	.prn(vcc));
defparam \prev_logical_channel[0] .is_wysiwyg = "true";
defparam \prev_logical_channel[0] .power_up = "low";

dffeas \prev_logical_channel[1] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[1]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[1]~q ),
	.prn(vcc));
defparam \prev_logical_channel[1] .is_wysiwyg = "true";
defparam \prev_logical_channel[1] .power_up = "low";

dffeas \prev_logical_channel[2] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[2]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[2]~q ),
	.prn(vcc));
defparam \prev_logical_channel[2] .is_wysiwyg = "true";
defparam \prev_logical_channel[2] .power_up = "low";

cyclonev_lcell_comb \Equal2~2 (
	.dataa(!\prev_logical_channel[0]~q ),
	.datab(!\alt_cal_inst|alt_cal_channel[0]~q ),
	.datac(!\prev_logical_channel[1]~q ),
	.datad(!\alt_cal_inst|alt_cal_channel[1]~q ),
	.datae(!\prev_logical_channel[2]~q ),
	.dataf(!\alt_cal_inst|alt_cal_channel[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~2 .extended_lut = "off";
defparam \Equal2~2 .lut_mask = 64'h9009000000009009;
defparam \Equal2~2 .shared_arith = "off";

dffeas \prev_logical_channel[3] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[3]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[3]~q ),
	.prn(vcc));
defparam \prev_logical_channel[3] .is_wysiwyg = "true";
defparam \prev_logical_channel[3] .power_up = "low";

dffeas \prev_logical_channel[4] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[4]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[4]~q ),
	.prn(vcc));
defparam \prev_logical_channel[4] .is_wysiwyg = "true";
defparam \prev_logical_channel[4] .power_up = "low";

dffeas \prev_logical_channel[5] (
	.clk(mgmt_clk_clk),
	.d(\alt_cal_inst|alt_cal_channel[5]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector0~3_combout ),
	.q(\prev_logical_channel[5]~q ),
	.prn(vcc));
defparam \prev_logical_channel[5] .is_wysiwyg = "true";
defparam \prev_logical_channel[5] .power_up = "low";

cyclonev_lcell_comb \Equal2~3 (
	.dataa(!\prev_logical_channel[3]~q ),
	.datab(!\alt_cal_inst|alt_cal_channel[3]~q ),
	.datac(!\prev_logical_channel[4]~q ),
	.datad(!\alt_cal_inst|alt_cal_channel[4]~q ),
	.datae(!\prev_logical_channel[5]~q ),
	.dataf(!\alt_cal_inst|alt_cal_channel[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~3 .extended_lut = "off";
defparam \Equal2~3 .lut_mask = 64'h9009000000009009;
defparam \Equal2~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~7 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\always1~0_combout ),
	.datac(!\Equal2~0_combout ),
	.datad(!\Equal2~1_combout ),
	.datae(!\Equal2~2_combout ),
	.dataf(!\Equal2~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~7 .extended_lut = "off";
defparam \Selector45~7 .lut_mask = 64'h1111111111111151;
defparam \Selector45~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.RELEASE_PMUTEX_STATE~q ),
	.datac(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datad(!\Selector45~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h2F222F222F222F22;
defparam \Selector28~0 .shared_arith = "off";

dffeas \state.RELEASE_PMUTEX_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.RELEASE_PMUTEX_STATE~q ),
	.prn(vcc));
defparam \state.RELEASE_PMUTEX_STATE .is_wysiwyg = "true";
defparam \state.RELEASE_PMUTEX_STATE .power_up = "low";

dffeas \state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.RELEASE_PMUTEX_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.prn(vcc));
defparam \state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE .is_wysiwyg = "true";
defparam \state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE .power_up = "low";

dffeas \state.RELEASE_PHY_RESET_OVERRIDE_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.RELEASE_PHY_RESET_OVERRIDE_DATA_STATE~q ),
	.prn(vcc));
defparam \state.RELEASE_PHY_RESET_OVERRIDE_DATA_STATE .is_wysiwyg = "true";
defparam \state.RELEASE_PHY_RESET_OVERRIDE_DATA_STATE .power_up = "low";

dffeas \state.RELEASE_PHY_RESET_OVERRIDE_START_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.RELEASE_PHY_RESET_OVERRIDE_DATA_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.RELEASE_PHY_RESET_OVERRIDE_START_STATE~q ),
	.prn(vcc));
defparam \state.RELEASE_PHY_RESET_OVERRIDE_START_STATE .is_wysiwyg = "true";
defparam \state.RELEASE_PHY_RESET_OVERRIDE_START_STATE .power_up = "low";

dffeas \state.RELEASE_OC_CALEN_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.RELEASE_PHY_RESET_OVERRIDE_START_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.RELEASE_OC_CALEN_DATA_STATE~q ),
	.prn(vcc));
defparam \state.RELEASE_OC_CALEN_DATA_STATE .is_wysiwyg = "true";
defparam \state.RELEASE_OC_CALEN_DATA_STATE .power_up = "low";

dffeas \state.RELEASE_OC_CALEN_START_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.RELEASE_OC_CALEN_DATA_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.RELEASE_OC_CALEN_START_STATE~q ),
	.prn(vcc));
defparam \state.RELEASE_OC_CALEN_START_STATE .is_wysiwyg = "true";
defparam \state.RELEASE_OC_CALEN_START_STATE .power_up = "low";

dffeas \state.RELEASE_OC_CALEN_DONE_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.RELEASE_OC_CALEN_START_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.RELEASE_OC_CALEN_DONE_STATE~q ),
	.prn(vcc));
defparam \state.RELEASE_OC_CALEN_DONE_STATE .is_wysiwyg = "true";
defparam \state.RELEASE_OC_CALEN_DONE_STATE .power_up = "low";

cyclonev_lcell_comb \Selector15~0 (
	.dataa(!basic_reconfig_readdata_2),
	.datab(!Equal8),
	.datac(!\state.CHECK_PHY_ADDR_STATE~q ),
	.datad(!\state.CHECK_REQ_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "off";
defparam \Selector15~0 .lut_mask = 64'h03AB03AB03AB03AB;
defparam \Selector15~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~1 (
	.dataa(!\state.000000~q ),
	.datab(!\always1~0_combout ),
	.datac(!\master_write~0_combout ),
	.datad(!\state.RELEASE_OC_CALEN_DONE_STATE~q ),
	.datae(!\Selector15~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~1 .extended_lut = "off";
defparam \Selector15~1 .lut_mask = 64'hDDD00000DDD00000;
defparam \Selector15~1 .shared_arith = "off";

dffeas \state.000000 (
	.clk(mgmt_clk_clk),
	.d(\Selector15~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.000000~q ),
	.prn(vcc));
defparam \state.000000 .is_wysiwyg = "true";
defparam \state.000000 .power_up = "low";

cyclonev_lcell_comb \Selector16~1 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal2~1_combout ),
	.datac(!\Equal2~2_combout ),
	.datad(!\Equal2~3_combout ),
	.datae(!\Selector16~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~1 .extended_lut = "off";
defparam \Selector16~1 .lut_mask = 64'h0000000200000002;
defparam \Selector16~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~2 (
	.dataa(!\state.000000~q ),
	.datab(!\always1~0_combout ),
	.datac(!\master_write~0_combout ),
	.datad(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datae(!\Selector16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~2 .extended_lut = "off";
defparam \Selector16~2 .lut_mask = 64'h88F8CCFC88F8CCFC;
defparam \Selector16~2 .shared_arith = "off";

dffeas \state.LOGICAL_ADDRESS_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector16~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOGICAL_ADDRESS_STATE~q ),
	.prn(vcc));
defparam \state.LOGICAL_ADDRESS_STATE .is_wysiwyg = "true";
defparam \state.LOGICAL_ADDRESS_STATE .power_up = "low";

dffeas \state.READ_PHY_ADDR_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.LOGICAL_ADDRESS_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.READ_PHY_ADDR_STATE~q ),
	.prn(vcc));
defparam \state.READ_PHY_ADDR_STATE .is_wysiwyg = "true";
defparam \state.READ_PHY_ADDR_STATE .power_up = "low";

cyclonev_lcell_comb \state~44 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.READ_PHY_ADDR_STATE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~44 .extended_lut = "off";
defparam \state~44 .lut_mask = 64'h1111111111111111;
defparam \state~44 .shared_arith = "off";

dffeas \state.CHECK_PHY_ADDR_STATE (
	.clk(mgmt_clk_clk),
	.d(\state~44_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CHECK_PHY_ADDR_STATE~q ),
	.prn(vcc));
defparam \state.CHECK_PHY_ADDR_STATE .is_wysiwyg = "true";
defparam \state.CHECK_PHY_ADDR_STATE .power_up = "low";

cyclonev_lcell_comb \Selector21~0 (
	.dataa(!Equal8),
	.datab(!\state.CHECK_PHY_ADDR_STATE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~0 .extended_lut = "off";
defparam \Selector21~0 .lut_mask = 64'h2222222222222222;
defparam \Selector21~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector21~1 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.datac(!\Selector21~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~1 .extended_lut = "off";
defparam \Selector21~1 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \Selector21~1 .shared_arith = "off";

dffeas \state.SET_ADDR_OFFSET_REQ_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector21~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.prn(vcc));
defparam \state.SET_ADDR_OFFSET_REQ_STATE .is_wysiwyg = "true";
defparam \state.SET_ADDR_OFFSET_REQ_STATE .power_up = "low";

dffeas \state.REQUEST_CONTROL_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.REQUEST_CONTROL_STATE~q ),
	.prn(vcc));
defparam \state.REQUEST_CONTROL_STATE .is_wysiwyg = "true";
defparam \state.REQUEST_CONTROL_STATE .power_up = "low";

cyclonev_lcell_comb \Selector23~0 (
	.dataa(!master_read1),
	.datab(!\master_write~0_combout ),
	.datac(!\state.REQUEST_CONTROL_STATE~q ),
	.datad(!\state.READ_REQ_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h03EF03EF03EF03EF;
defparam \Selector23~0 .shared_arith = "off";

dffeas \state.READ_REQ_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READ_REQ_DATA_STATE~q ),
	.prn(vcc));
defparam \state.READ_REQ_DATA_STATE .is_wysiwyg = "true";
defparam \state.READ_REQ_DATA_STATE .power_up = "low";

cyclonev_lcell_comb \state~45 (
	.dataa(!master_read1),
	.datab(!\master_write~0_combout ),
	.datac(!\state.READ_REQ_DATA_STATE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~45 .extended_lut = "off";
defparam \state~45 .lut_mask = 64'h0101010101010101;
defparam \state~45 .shared_arith = "off";

dffeas \state.CHECK_REQ_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\state~45_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CHECK_REQ_DATA_STATE~q ),
	.prn(vcc));
defparam \state.CHECK_REQ_DATA_STATE .is_wysiwyg = "true";
defparam \state.CHECK_REQ_DATA_STATE .power_up = "low";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!basic_reconfig_readdata_2),
	.datac(!\state.CHECK_PMUTEX_STATE~q ),
	.datad(!\state.CHECK_REQ_DATA_STATE~q ),
	.datae(!\pmutex_acquired~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'h0A3B0A0A0A3B0A0A;
defparam \Selector26~0 .shared_arith = "off";

dffeas \state.ACQUIRE_PMUTEX_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector26~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ACQUIRE_PMUTEX_STATE~q ),
	.prn(vcc));
defparam \state.ACQUIRE_PMUTEX_STATE .is_wysiwyg = "true";
defparam \state.ACQUIRE_PMUTEX_STATE .power_up = "low";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!master_read1),
	.datab(!\state.ACQUIRE_PMUTEX_STATE~q ),
	.datac(!\master_write~0_combout ),
	.datad(!\state.READ_PMUTEX_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h33FB33FB33FB33FB;
defparam \Selector27~0 .shared_arith = "off";

dffeas \state.READ_PMUTEX_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector27~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READ_PMUTEX_STATE~q ),
	.prn(vcc));
defparam \state.READ_PMUTEX_STATE .is_wysiwyg = "true";
defparam \state.READ_PMUTEX_STATE .power_up = "low";

cyclonev_lcell_comb \state~43 (
	.dataa(!master_read1),
	.datab(!\master_write~0_combout ),
	.datac(!\state.READ_PMUTEX_STATE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~43 .extended_lut = "off";
defparam \state~43 .lut_mask = 64'h0101010101010101;
defparam \state~43 .shared_arith = "off";

dffeas \state.CHECK_PMUTEX_STATE (
	.clk(mgmt_clk_clk),
	.d(\state~43_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CHECK_PMUTEX_STATE~q ),
	.prn(vcc));
defparam \state.CHECK_PMUTEX_STATE .is_wysiwyg = "true";
defparam \state.CHECK_PMUTEX_STATE .power_up = "low";

cyclonev_lcell_comb \Selector38~0 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!\state.CHECK_PMUTEX_STATE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~0 .extended_lut = "off";
defparam \Selector38~0 .lut_mask = 64'h1111111111111111;
defparam \Selector38~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector38~1 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datac(!\Selector38~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~1 .extended_lut = "off";
defparam \Selector38~1 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \Selector38~1 .shared_arith = "off";

dffeas \state.SET_PHY_RESET_OVERRIDE_ADDR_STATE (
	.clk(mgmt_clk_clk),
	.d(\Selector38~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.prn(vcc));
defparam \state.SET_PHY_RESET_OVERRIDE_ADDR_STATE .is_wysiwyg = "true";
defparam \state.SET_PHY_RESET_OVERRIDE_ADDR_STATE .power_up = "low";

dffeas \state.SET_PHY_RESET_OVERRIDE_DATA_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.SET_PHY_RESET_OVERRIDE_DATA_STATE~q ),
	.prn(vcc));
defparam \state.SET_PHY_RESET_OVERRIDE_DATA_STATE .is_wysiwyg = "true";
defparam \state.SET_PHY_RESET_OVERRIDE_DATA_STATE .power_up = "low";

dffeas \state.SET_PHY_RESET_OVERRIDE_START_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.SET_PHY_RESET_OVERRIDE_DATA_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.SET_PHY_RESET_OVERRIDE_START_STATE~q ),
	.prn(vcc));
defparam \state.SET_PHY_RESET_OVERRIDE_START_STATE .is_wysiwyg = "true";
defparam \state.SET_PHY_RESET_OVERRIDE_START_STATE .power_up = "low";

dffeas \state.GET_TESTBUS_ADDR_STATE (
	.clk(mgmt_clk_clk),
	.d(\state.SET_PHY_RESET_OVERRIDE_START_STATE~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\master_write~0_combout ),
	.q(\state.GET_TESTBUS_ADDR_STATE~q ),
	.prn(vcc));
defparam \state.GET_TESTBUS_ADDR_STATE .is_wysiwyg = "true";
defparam \state.GET_TESTBUS_ADDR_STATE .power_up = "low";

cyclonev_lcell_comb \Selector78~0 (
	.dataa(!\state.CONTROL_STATE~q ),
	.datab(!\state.START_OC_CALEN_STATE~q ),
	.datac(!\state.RELEASE_OC_CALEN_START_STATE~q ),
	.datad(!\state.SET_PHY_RESET_OVERRIDE_DATA_STATE~q ),
	.datae(!\state.RELEASE_PHY_RESET_OVERRIDE_DATA_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~0 .extended_lut = "off";
defparam \Selector78~0 .lut_mask = 64'h8000000080000000;
defparam \Selector78~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\state.SET_OC_CALEN_DATA_STATE~q ),
	.datab(!\state.RELEASE_OC_CALEN_DATA_STATE~q ),
	.datac(!\state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h8080808080808080;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!\state.SET_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datab(!\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.datac(!\state.SET_OC_CALEN_ADDR_STATE~q ),
	.datad(!\state.RELEASE_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h8000800080008000;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!\state.REQUEST_CONTROL_STATE~q ),
	.datab(!\state.GET_TESTBUS_DATA_STATE~q ),
	.datac(!\Selector78~0_combout ),
	.datad(!\Selector1~0_combout ),
	.datae(!\Selector1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h0000000800000008;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datab(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datac(!\Selector1~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h0808080808080808;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\Selector1~3_combout ),
	.datab(!\state.RELEASE_PMUTEX_STATE~q ),
	.datac(!\state.WRITE_DATA_STATE~q ),
	.datad(!\state.ADDRESS_OFFSET_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h4000400040004000;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~1 (
	.dataa(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datab(!\state.READ_DATA_STATE~q ),
	.datac(!\state.BUSY_STATE~q ),
	.datad(!\state.READ_PHY_ADDR_STATE~q ),
	.datae(!\state.RELEASE_OC_CALEN_DONE_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~1 .extended_lut = "off";
defparam \Selector0~1 .lut_mask = 64'h8000000080000000;
defparam \Selector0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~2 (
	.dataa(!master_read1),
	.datab(!\master_write~0_combout ),
	.datac(!\Selector0~1_combout ),
	.datad(!\state.READ_REQ_DATA_STATE~q ),
	.datae(!\state.READ_PMUTEX_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~2 .extended_lut = "off";
defparam \Selector0~2 .lut_mask = 64'h3F2222223F222222;
defparam \Selector0~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~4 (
	.dataa(!master_write1),
	.datab(!\alt_cal_inst|alt_cal_busy~q ),
	.datac(!\alt_cal_inst|write_reg~q ),
	.datad(!\alt_cal_inst|read~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~4 .extended_lut = "off";
defparam \Selector0~4 .lut_mask = 64'h2000200020002000;
defparam \Selector0~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~5 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!master_write1),
	.datac(!\state.CHECK_PMUTEX_STATE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~5 .extended_lut = "off";
defparam \Selector0~5 .lut_mask = 64'h0707070707070707;
defparam \Selector0~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~6 (
	.dataa(!\state.ACQUIRE_PMUTEX_STATE~q ),
	.datab(!\Selector0~3_combout ),
	.datac(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datad(!\Selector0~4_combout ),
	.datae(!\Selector0~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~6 .extended_lut = "off";
defparam \Selector0~6 .lut_mask = 64'h8088000080880000;
defparam \Selector0~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~7 (
	.dataa(!master_write1),
	.datab(!\master_write~0_combout ),
	.datac(!\Selector0~0_combout ),
	.datad(!\Selector0~2_combout ),
	.datae(!\Selector0~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~7 .extended_lut = "off";
defparam \Selector0~7 .lut_mask = 64'hFFFF7570FFFF7570;
defparam \Selector0~7 .shared_arith = "off";

cyclonev_lcell_comb \offset_cancellation_done~2 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.000000~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_cancellation_done~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_cancellation_done~2 .extended_lut = "off";
defparam \offset_cancellation_done~2 .lut_mask = 64'h7777777777777777;
defparam \offset_cancellation_done~2 .shared_arith = "off";

cyclonev_lcell_comb \master_address~0 (
	.dataa(!master_write1),
	.datab(!master_read1),
	.datac(!\master_write~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_address~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_address~0 .extended_lut = "off";
defparam \master_address~0 .lut_mask = 64'h0404040404040404;
defparam \master_address~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~0 (
	.dataa(!\state.REQUEST_CONTROL_STATE~q ),
	.datab(!\state.GET_TESTBUS_DATA_STATE~q ),
	.datac(!\Selector78~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~0 .extended_lut = "off";
defparam \Selector45~0 .lut_mask = 64'h0808080808080808;
defparam \Selector45~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector44~0 (
	.dataa(!\master_write~0_combout ),
	.datab(!\Selector45~0_combout ),
	.datac(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datad(!\state.READ_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector44~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector44~0 .extended_lut = "off";
defparam \Selector44~0 .lut_mask = 64'h8AAA8AAA8AAA8AAA;
defparam \Selector44~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr2~0 (
	.dataa(!\state.CHECK_PHY_ADDR_STATE~q ),
	.datab(!\state.CHECK_REQ_DATA_STATE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr2~0 .extended_lut = "off";
defparam \WideOr2~0 .lut_mask = 64'h7777777777777777;
defparam \WideOr2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector44~1 (
	.dataa(!\state.BUSY_STATE~q ),
	.datab(!\state.READ_PHY_ADDR_STATE~q ),
	.datac(!\state.RELEASE_OC_CALEN_DONE_STATE~q ),
	.datad(!\state.READ_REQ_DATA_STATE~q ),
	.datae(!\WideOr2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector44~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector44~1 .extended_lut = "off";
defparam \Selector44~1 .lut_mask = 64'h8000000080000000;
defparam \Selector44~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector44~2 (
	.dataa(!\always1~0_combout ),
	.datab(!\state.CHECK_PMUTEX_STATE~q ),
	.datac(!\Selector44~0_combout ),
	.datad(!\Selector14~0_combout ),
	.datae(!\Selector44~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector44~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector44~2 .extended_lut = "off";
defparam \Selector44~2 .lut_mask = 64'h000080C0000080C0;
defparam \Selector44~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~1 (
	.dataa(!\state.SET_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datab(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datac(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datad(!\state.WRITE_DATA_STATE~q ),
	.datae(!\state.ADDRESS_OFFSET_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~1 .extended_lut = "off";
defparam \Selector45~1 .lut_mask = 64'h8000000080000000;
defparam \Selector45~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~2 (
	.dataa(!\state.SET_OC_CALEN_ADDR_STATE~q ),
	.datab(!\state.RELEASE_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datac(!\state.RELEASE_OC_CALEN_DATA_STATE~q ),
	.datad(!\state.RELEASE_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datae(!\Selector45~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~2 .extended_lut = "off";
defparam \Selector45~2 .lut_mask = 64'h0000800000008000;
defparam \Selector45~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~3 (
	.dataa(!\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.datab(!\state.SET_OC_CALEN_DATA_STATE~q ),
	.datac(!\Selector45~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~3 .extended_lut = "off";
defparam \Selector45~3 .lut_mask = 64'h0808080808080808;
defparam \Selector45~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector44~4 (
	.dataa(!\Selector45~3_combout ),
	.datab(!\state.RELEASE_PMUTEX_STATE~q ),
	.datac(!\state.BUSY_STATE~q ),
	.datad(!\Selector38~0_combout ),
	.datae(!\master_write~0_combout ),
	.dataf(!\write_read_control~q ),
	.datag(!master_address_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector44~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector44~4 .extended_lut = "on";
defparam \Selector44~4 .lut_mask = 64'h0BFFBFFF0BFFBBFF;
defparam \Selector44~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector44~3 (
	.dataa(!master_address_2),
	.datab(!\state.READ_REQ_DATA_STATE~q ),
	.datac(!\state.READ_PMUTEX_STATE~q ),
	.datad(!\master_address~0_combout ),
	.datae(!\Selector44~2_combout ),
	.dataf(!\Selector44~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector44~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector44~3 .extended_lut = "off";
defparam \Selector44~3 .lut_mask = 64'h55770533FFFFFFFF;
defparam \Selector44~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector46~0 (
	.dataa(!\Selector45~0_combout ),
	.datab(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datac(!\Selector1~0_combout ),
	.datad(!\state.WRITE_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~0 .extended_lut = "off";
defparam \Selector46~0 .lut_mask = 64'h0400040004000400;
defparam \Selector46~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~4 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!\state.CHECK_PMUTEX_STATE~q ),
	.datac(!\state.READ_PHY_ADDR_STATE~q ),
	.datad(!\state.RELEASE_OC_CALEN_DONE_STATE~q ),
	.datae(!\state.READ_PMUTEX_STATE~q ),
	.dataf(!\WideOr2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~4 .extended_lut = "off";
defparam \Selector45~4 .lut_mask = 64'hD000000000000000;
defparam \Selector45~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector46~1 (
	.dataa(!\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.datab(!\state.SET_OC_CALEN_ADDR_STATE~q ),
	.datac(!\state.RELEASE_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datad(!\state.RELEASE_PMUTEX_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~1 .extended_lut = "off";
defparam \Selector46~1 .lut_mask = 64'h8000800080008000;
defparam \Selector46~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector46~2 (
	.dataa(!\state.SET_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datab(!\state.ADDRESS_OFFSET_STATE~q ),
	.datac(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datad(!\state.READ_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~2 .extended_lut = "off";
defparam \Selector46~2 .lut_mask = 64'h8000800080008000;
defparam \Selector46~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector46~3 (
	.dataa(!\state.000000~q ),
	.datab(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datac(!\state.BUSY_STATE~q ),
	.datad(!\state.READ_REQ_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~3 .extended_lut = "off";
defparam \Selector46~3 .lut_mask = 64'h4000400040004000;
defparam \Selector46~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector46~4 (
	.dataa(!\master_write~0_combout ),
	.datab(!\Selector45~4_combout ),
	.datac(!\Selector46~1_combout ),
	.datad(!\Selector46~2_combout ),
	.datae(!\Selector46~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~4 .extended_lut = "off";
defparam \Selector46~4 .lut_mask = 64'hFFFFEEECFFFFEEEC;
defparam \Selector46~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector46~5 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.000000~q ),
	.datac(!\state.ACQUIRE_PMUTEX_STATE~q ),
	.datad(!\always1~0_combout ),
	.datae(!\state.WAIT_FOR_NEXT_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~5 .extended_lut = "off";
defparam \Selector46~5 .lut_mask = 64'hCF0FFFAFCF0FFFAF;
defparam \Selector46~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~4 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.BUSY_STATE~q ),
	.datac(!\state.READ_REQ_DATA_STATE~q ),
	.datad(!\state.READ_PMUTEX_STATE~q ),
	.datae(!\master_address~0_combout ),
	.dataf(!\write_read_control~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~4 .extended_lut = "off";
defparam \Selector1~4 .lut_mask = 64'hEEEEE000FFFFF000;
defparam \Selector1~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector46~6 (
	.dataa(!\Selector46~0_combout ),
	.datab(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datac(!\Selector46~4_combout ),
	.datad(!\Selector46~5_combout ),
	.datae(!master_address_0),
	.dataf(!\Selector1~4_combout ),
	.datag(!\master_write~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~6 .extended_lut = "on";
defparam \Selector46~6 .lut_mask = 64'hFFFFFFFF0BFFBFFF;
defparam \Selector46~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~5 (
	.dataa(!\state.000000~q ),
	.datab(!\alt_cal_inst|write_reg~q ),
	.datac(!\alt_cal_inst|read~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\Selector45~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~5 .extended_lut = "off";
defparam \Selector45~5 .lut_mask = 64'h00007F3F00007F3F;
defparam \Selector45~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~6 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.BUSY_STATE~q ),
	.datac(!\state.READ_REQ_DATA_STATE~q ),
	.datad(!\master_address~0_combout ),
	.datae(!\write_read_control~q ),
	.dataf(!\Selector45~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~6 .extended_lut = "off";
defparam \Selector45~6 .lut_mask = 64'h00000000D0DDC0CC;
defparam \Selector45~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~8 (
	.dataa(!\state.RELEASE_PMUTEX_STATE~q ),
	.datab(!\state.READ_DATA_STATE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~8 .extended_lut = "off";
defparam \Selector45~8 .lut_mask = 64'h8888888888888888;
defparam \Selector45~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~9 (
	.dataa(!master_address_1),
	.datab(!\master_write~0_combout ),
	.datac(!\Selector45~8_combout ),
	.datad(!\Selector45~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~9 .extended_lut = "off";
defparam \Selector45~9 .lut_mask = 64'h4440444044404440;
defparam \Selector45~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~10 (
	.dataa(!\state.ACQUIRE_PMUTEX_STATE~q ),
	.datab(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datac(!\state.READ_PMUTEX_STATE~q ),
	.datad(!\master_address~0_combout ),
	.datae(!\Selector45~7_combout ),
	.dataf(!\Selector45~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~10 .extended_lut = "off";
defparam \Selector45~10 .lut_mask = 64'h8880AAA000000000;
defparam \Selector45~10 .shared_arith = "off";

cyclonev_lcell_comb \Selector45~11 (
	.dataa(!master_address_1),
	.datab(!\master_write~0_combout ),
	.datac(!\Selector45~0_combout ),
	.datad(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datae(!\Selector45~6_combout ),
	.dataf(!\Selector45~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~11 .extended_lut = "off";
defparam \Selector45~11 .lut_mask = 64'hFFFFFFFF75777077;
defparam \Selector45~11 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~5 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~5 .extended_lut = "off";
defparam \Selector1~5 .lut_mask = 64'h1111111111111111;
defparam \Selector1~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~6 (
	.dataa(!\always1~0_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\Equal2~1_combout ),
	.datad(!\Equal2~2_combout ),
	.datae(!\Equal2~3_combout ),
	.dataf(!\Selector16~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~6 .extended_lut = "off";
defparam \Selector1~6 .lut_mask = 64'h000000005555555D;
defparam \Selector1~6 .shared_arith = "off";

cyclonev_lcell_comb \WideOr34~0 (
	.dataa(!\state.BUSY_STATE~q ),
	.datab(!\state.READ_PHY_ADDR_STATE~q ),
	.datac(!\state.RELEASE_OC_CALEN_DONE_STATE~q ),
	.datad(!\state.READ_REQ_DATA_STATE~q ),
	.datae(!\state.READ_PMUTEX_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr34~0 .extended_lut = "off";
defparam \WideOr34~0 .lut_mask = 64'h8000000080000000;
defparam \WideOr34~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~7 (
	.dataa(!\state.RELEASE_PMUTEX_STATE~q ),
	.datab(!\state.WRITE_DATA_STATE~q ),
	.datac(!\state.ADDRESS_OFFSET_STATE~q ),
	.datad(!\state.READ_DATA_STATE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~7 .extended_lut = "off";
defparam \Selector1~7 .lut_mask = 64'h8000800080008000;
defparam \Selector1~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~8 (
	.dataa(!\master_write~0_combout ),
	.datab(!\Selector1~3_combout ),
	.datac(!\WideOr34~0_combout ),
	.datad(!\Selector1~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~8 .extended_lut = "off";
defparam \Selector1~8 .lut_mask = 64'hAAA8AAA8AAA8AAA8;
defparam \Selector1~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~9 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!\state.CHECK_PMUTEX_STATE~q ),
	.datac(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~9 .extended_lut = "off";
defparam \Selector1~9 .lut_mask = 64'hD0D0D0D0D0D0D0D0;
defparam \Selector1~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~10 (
	.dataa(!master_read1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector1~5_combout ),
	.datad(!\Selector1~6_combout ),
	.datae(!\Selector1~8_combout ),
	.dataf(!\Selector1~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~10 .extended_lut = "off";
defparam \Selector1~10 .lut_mask = 64'hDFDFDFDFCFDFDFDF;
defparam \Selector1~10 .shared_arith = "off";

cyclonev_lcell_comb \oc_started~0 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\oc_started~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oc_started~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oc_started~0 .extended_lut = "off";
defparam \oc_started~0 .lut_mask = 64'h7777777777777777;
defparam \oc_started~0 .shared_arith = "off";

dffeas oc_started(
	.clk(mgmt_clk_clk),
	.d(\oc_started~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\oc_started~q ),
	.prn(vcc));
defparam oc_started.is_wysiwyg = "true";
defparam oc_started.power_up = "low";

cyclonev_lcell_comb WideOr34(
	.dataa(!\state.LOGICAL_ADDRESS_STATE~q ),
	.datab(!\WideOr2~0_combout ),
	.datac(!\WideOr34~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr34~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr34.extended_lut = "off";
defparam WideOr34.lut_mask = 64'h0808080808080808;
defparam WideOr34.shared_arith = "off";

cyclonev_lcell_comb \Selector67~0 (
	.dataa(!\always1~0_combout ),
	.datab(!\state.CHECK_PMUTEX_STATE~q ),
	.datac(!\Selector14~0_combout ),
	.datad(!\WideOr34~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector67~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector67~0 .extended_lut = "off";
defparam \Selector67~0 .lut_mask = 64'h008C008C008C008C;
defparam \Selector67~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector77~0 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_OC_CALEN_ADDR_STATE~q ),
	.datac(!\state.RELEASE_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datad(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datae(!\state.RELEASE_PMUTEX_STATE~q ),
	.dataf(!master_write_data_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector77~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector77~0 .extended_lut = "off";
defparam \Selector77~0 .lut_mask = 64'hEAAAAAAAC0000000;
defparam \Selector77~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector77~1 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.WRITE_DATA_STATE~q ),
	.datac(!\state.ADDRESS_OFFSET_STATE~q ),
	.datad(!\alt_cal_inst|address[1]~q ),
	.datae(!\alt_cal_inst|dataout[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector77~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector77~1 .extended_lut = "off";
defparam \Selector77~1 .lut_mask = 64'h0005111500051115;
defparam \Selector77~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector77~2 (
	.dataa(!\state.SET_PHY_RESET_OVERRIDE_START_STATE~q ),
	.datab(!\state.ADDRESS_OFFSET_STATE~q ),
	.datac(!\state.READ_DATA_STATE~q ),
	.datad(!\Selector46~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector77~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector77~2 .extended_lut = "off";
defparam \Selector77~2 .lut_mask = 64'h0080008000800080;
defparam \Selector77~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector77~3 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.datac(!\Selector77~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector77~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector77~3 .extended_lut = "off";
defparam \Selector77~3 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \Selector77~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector77~4 (
	.dataa(!\state.000000~q ),
	.datab(!\always1~0_combout ),
	.datac(!\alt_cal_inst|alt_cal_channel[1]~q ),
	.datad(!\Selector38~0_combout ),
	.datae(!\Selector16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector77~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector77~4 .extended_lut = "off";
defparam \Selector77~4 .lut_mask = 64'hF700F300F700F300;
defparam \Selector77~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector77~5 (
	.dataa(!master_write_data_1),
	.datab(!\Selector67~0_combout ),
	.datac(!\Selector77~0_combout ),
	.datad(!\Selector77~1_combout ),
	.datae(!\Selector77~3_combout ),
	.dataf(!\Selector77~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector77~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector77~5 .extended_lut = "off";
defparam \Selector77~5 .lut_mask = 64'hFFFFFFFFF4FFF5FF;
defparam \Selector77~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector76~0 (
	.dataa(!\state.000000~q ),
	.datab(!\always1~0_combout ),
	.datac(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datad(!\alt_cal_inst|alt_cal_channel[2]~q ),
	.datae(!master_write_data_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~0 .extended_lut = "off";
defparam \Selector76~0 .lut_mask = 64'h008C23AF008C23AF;
defparam \Selector76~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector76~1 (
	.dataa(!\state.WRITE_DATA_STATE~q ),
	.datab(!\state.ADDRESS_OFFSET_STATE~q ),
	.datac(!\alt_cal_inst|address[1]~q ),
	.datad(!\alt_cal_inst|dataout[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~1 .extended_lut = "off";
defparam \Selector76~1 .lut_mask = 64'h0357035703570357;
defparam \Selector76~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector76~2 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datac(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datad(!\Selector76~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~2 .extended_lut = "off";
defparam \Selector76~2 .lut_mask = 64'h1555155515551555;
defparam \Selector76~2 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[7]~0 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!\state.CHECK_PMUTEX_STATE~q ),
	.datac(!\WideOr34~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[7]~0 .extended_lut = "off";
defparam \master_write_data[7]~0 .lut_mask = 64'h0D0D0D0D0D0D0D0D;
defparam \master_write_data[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector76~3 (
	.dataa(!\Selector1~2_combout ),
	.datab(!\Selector1~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~3 .extended_lut = "off";
defparam \Selector76~3 .lut_mask = 64'h1111111111111111;
defparam \Selector76~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector76~4 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datac(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datad(!master_write_data_2),
	.datae(!\master_write_data[7]~0_combout ),
	.dataf(!\Selector76~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~4 .extended_lut = "off";
defparam \Selector76~4 .lut_mask = 64'h00FF00BF00FF003F;
defparam \Selector76~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector76~5 (
	.dataa(!\state.ACQUIRE_PMUTEX_STATE~q ),
	.datab(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datac(!\Selector45~7_combout ),
	.datad(!\Selector76~0_combout ),
	.datae(!\Selector76~2_combout ),
	.dataf(!\Selector76~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~5 .extended_lut = "off";
defparam \Selector76~5 .lut_mask = 64'h75FFFFFFFFFFFFFF;
defparam \Selector76~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector78~1 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.CONTROL_STATE~q ),
	.datac(!\write_read_control~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~1 .extended_lut = "off";
defparam \Selector78~1 .lut_mask = 64'h1010101010101010;
defparam \Selector78~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector78~2 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.datac(!\state.SET_OC_CALEN_DATA_STATE~q ),
	.datad(!\state.REQUEST_CONTROL_STATE~q ),
	.datae(!master_write_data_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~2 .extended_lut = "off";
defparam \Selector78~2 .lut_mask = 64'hEAAAC000EAAAC000;
defparam \Selector78~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector78~3 (
	.dataa(!\state.WRITE_DATA_STATE~q ),
	.datab(!\state.ADDRESS_OFFSET_STATE~q ),
	.datac(!\alt_cal_inst|dataout[0]~q ),
	.datad(!\alt_cal_inst|address[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~3 .extended_lut = "off";
defparam \Selector78~3 .lut_mask = 64'h0537053705370537;
defparam \Selector78~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector78~4 (
	.dataa(!\state.GET_TESTBUS_DATA_STATE~q ),
	.datab(!\Selector78~0_combout ),
	.datac(!\Selector45~8_combout ),
	.datad(!\Selector45~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~4 .extended_lut = "off";
defparam \Selector78~4 .lut_mask = 64'h0002000200020002;
defparam \Selector78~4 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[7]~1 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.000000~q ),
	.datac(!\alt_cal_inst|write_reg~q ),
	.datad(!\alt_cal_inst|read~q ),
	.datae(!\state.WAIT_FOR_NEXT_STATE~q ),
	.dataf(!\master_write_data[7]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[7]~1 .extended_lut = "off";
defparam \master_write_data[7]~1 .lut_mask = 64'h000000003FFF2FFF;
defparam \master_write_data[7]~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector78~5 (
	.dataa(!\master_write~0_combout ),
	.datab(!master_write_data_0),
	.datac(!\Selector78~4_combout ),
	.datad(!\master_write_data[7]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~5 .extended_lut = "off";
defparam \Selector78~5 .lut_mask = 64'h3320332033203320;
defparam \Selector78~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector78~6 (
	.dataa(!\state.000000~q ),
	.datab(!\state.ACQUIRE_PMUTEX_STATE~q ),
	.datac(!\always1~0_combout ),
	.datad(!\alt_cal_inst|alt_cal_channel[0]~q ),
	.datae(!\Selector16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~6 .extended_lut = "off";
defparam \Selector78~6 .lut_mask = 64'hCC4CCC0CCC4CCC0C;
defparam \Selector78~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector78~7 (
	.dataa(!\master_write~0_combout ),
	.datab(!\Selector78~1_combout ),
	.datac(!\Selector78~2_combout ),
	.datad(!\Selector78~3_combout ),
	.datae(!\Selector78~5_combout ),
	.dataf(!\Selector78~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~7 .extended_lut = "off";
defparam \Selector78~7 .lut_mask = 64'hFFFFFFFFF3F7FFFF;
defparam \Selector78~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~0 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_ADDR_OFFSET_REQ_STATE~q ),
	.datac(!\state.GET_TESTBUS_DATA_STATE~q ),
	.datad(!\state.RELEASE_PMUTEX_STATE~q ),
	.datae(!master_write_data_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~0 .extended_lut = "off";
defparam \Selector75~0 .lut_mask = 64'hEAAAC000EAAAC000;
defparam \Selector75~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~1 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.WRITE_DATA_STATE~q ),
	.datac(!\state.ADDRESS_OFFSET_STATE~q ),
	.datad(!\alt_cal_inst|address[1]~q ),
	.datae(!\alt_cal_inst|dataout[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~1 .extended_lut = "off";
defparam \Selector75~1 .lut_mask = 64'h0005111500051115;
defparam \Selector75~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~2 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_OC_CALEN_DATA_STATE~q ),
	.datac(!\state.REQUEST_CONTROL_STATE~q ),
	.datad(!\Selector78~0_combout ),
	.datae(!\state.READ_DATA_STATE~q ),
	.dataf(!\Selector45~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~2 .extended_lut = "off";
defparam \Selector75~2 .lut_mask = 64'hAAAAAAAAAA2AAAAA;
defparam \Selector75~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~3 (
	.dataa(!\state.000000~q ),
	.datab(!\always1~0_combout ),
	.datac(!\alt_cal_inst|alt_cal_channel[3]~q ),
	.datad(!\Selector38~0_combout ),
	.datae(!\Selector16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~3 .extended_lut = "off";
defparam \Selector75~3 .lut_mask = 64'hF700F300F700F300;
defparam \Selector75~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~4 (
	.dataa(!master_write_data_3),
	.datab(!\Selector75~0_combout ),
	.datac(!\Selector75~1_combout ),
	.datad(!\Selector75~2_combout ),
	.datae(!\Selector67~0_combout ),
	.dataf(!\Selector75~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~4 .extended_lut = "off";
defparam \Selector75~4 .lut_mask = 64'hFFFFFFFFDFDFCFDF;
defparam \Selector75~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector74~0 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datac(!\state.WRITE_DATA_STATE~q ),
	.datad(!\state.ADDRESS_OFFSET_STATE~q ),
	.datae(!\alt_cal_inst|dataout[4]~q ),
	.dataf(!\alt_cal_inst|address[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector74~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector74~0 .extended_lut = "off";
defparam \Selector74~0 .lut_mask = 64'h1111151511551555;
defparam \Selector74~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector74~1 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datac(!\state.SET_PHY_RESET_OVERRIDE_ADDR_STATE~q ),
	.datad(!master_write_data_4),
	.datae(!\master_write_data[7]~1_combout ),
	.dataf(!\Selector76~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector74~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector74~1 .extended_lut = "off";
defparam \Selector74~1 .lut_mask = 64'h00FF00AF00FF002F;
defparam \Selector74~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector74~2 (
	.dataa(!\state.000000~q ),
	.datab(!\always1~0_combout ),
	.datac(!\alt_cal_inst|alt_cal_channel[4]~q ),
	.datad(!\Selector16~1_combout ),
	.datae(!\Selector74~0_combout ),
	.dataf(!\Selector74~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector74~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector74~2 .extended_lut = "off";
defparam \Selector74~2 .lut_mask = 64'h080CFFFFFFFFFFFF;
defparam \Selector74~2 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[7]~2 (
	.dataa(!\state.000000~q ),
	.datab(!\state.ACQUIRE_PMUTEX_STATE~q ),
	.datac(!\state.WRITE_DATA_STATE~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\state.WRITE_DONE_STATE~q ),
	.dataf(!\WideOr34~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[7]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[7]~2 .extended_lut = "off";
defparam \master_write_data[7]~2 .lut_mask = 64'h3333FFFF7333FFFF;
defparam \master_write_data[7]~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~4 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal2~1_combout ),
	.datac(!\Equal2~2_combout ),
	.datad(!\Equal2~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~4 .extended_lut = "off";
defparam \Equal2~4 .lut_mask = 64'h0002000200020002;
defparam \Equal2~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector73~0 (
	.dataa(!\master_write_data[7]~2_combout ),
	.datab(!\Equal2~4_combout ),
	.datac(!\alt_cal_inst|dataout[5]~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\state.WRITE_DATA_STATE~q ),
	.dataf(!\alt_cal_inst|alt_cal_busy~q ),
	.datag(!\alt_cal_inst|alt_cal_channel[5]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector73~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector73~0 .extended_lut = "on";
defparam \Selector73~0 .lut_mask = 64'h0A000A000A020A02;
defparam \Selector73~0 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[7]~3 (
	.dataa(!\Selector1~3_combout ),
	.datab(!\state.ADDRESS_OFFSET_STATE~q ),
	.datac(!\Selector45~8_combout ),
	.datad(!\Selector38~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[7]~3 .extended_lut = "off";
defparam \master_write_data[7]~3 .lut_mask = 64'hFB00FB00FB00FB00;
defparam \master_write_data[7]~3 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[7]~4 (
	.dataa(!mutex_grant),
	.datab(!basic_reconfig_waitrequest2),
	.datac(!\state.WRITE_DATA_STATE~q ),
	.datad(!\state.CHECK_PMUTEX_STATE~q ),
	.datae(!\master_write_data[7]~1_combout ),
	.dataf(!\master_write_data[7]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[7]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[7]~4 .extended_lut = "off";
defparam \master_write_data[7]~4 .lut_mask = 64'h0000F4F400004400;
defparam \master_write_data[7]~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector72~0 (
	.dataa(!\master_write_data[7]~2_combout ),
	.datab(!\Equal2~4_combout ),
	.datac(!\alt_cal_inst|dataout[6]~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\state.WRITE_DATA_STATE~q ),
	.dataf(!\alt_cal_inst|alt_cal_busy~q ),
	.datag(!\alt_cal_inst|alt_cal_channel[6]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector72~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector72~0 .extended_lut = "on";
defparam \Selector72~0 .lut_mask = 64'h0A000A000A020A02;
defparam \Selector72~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector71~0 (
	.dataa(!\master_write_data[7]~2_combout ),
	.datab(!\Equal2~4_combout ),
	.datac(!\alt_cal_inst|dataout[7]~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\state.WRITE_DATA_STATE~q ),
	.dataf(!\alt_cal_inst|alt_cal_busy~q ),
	.datag(!\alt_cal_inst|alt_cal_channel[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector71~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector71~0 .extended_lut = "on";
defparam \Selector71~0 .lut_mask = 64'h0A000A000A020A02;
defparam \Selector71~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector70~0 (
	.dataa(!\master_write_data[7]~2_combout ),
	.datab(!\Equal2~4_combout ),
	.datac(!\alt_cal_inst|dataout[8]~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\state.WRITE_DATA_STATE~q ),
	.dataf(!\alt_cal_inst|alt_cal_busy~q ),
	.datag(!\alt_cal_inst|alt_cal_channel[8]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector70~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector70~0 .extended_lut = "on";
defparam \Selector70~0 .lut_mask = 64'h0A000A000A020A02;
defparam \Selector70~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector69~0 (
	.dataa(!\master_write_data[7]~2_combout ),
	.datab(!\Equal2~4_combout ),
	.datac(!\alt_cal_inst|dataout[9]~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\state.WRITE_DATA_STATE~q ),
	.dataf(!\alt_cal_inst|alt_cal_busy~q ),
	.datag(!\alt_cal_inst|alt_cal_channel[9]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector69~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector69~0 .extended_lut = "on";
defparam \Selector69~0 .lut_mask = 64'h0A000A000A020A02;
defparam \Selector69~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector68~0 (
	.dataa(!\state.WRITE_DATA_STATE~q ),
	.datab(!\alt_cal_inst|dataout[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector68~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector68~0 .extended_lut = "off";
defparam \Selector68~0 .lut_mask = 64'h1111111111111111;
defparam \Selector68~0 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[15]~5 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\Selector1~3_combout ),
	.datae(!\state.ADDRESS_OFFSET_STATE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[15]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[15]~5 .extended_lut = "off";
defparam \master_write_data[15]~5 .lut_mask = 64'h0400040404000404;
defparam \master_write_data[15]~5 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[15]~7 (
	.dataa(!\state.000000~q ),
	.datab(!\alt_cal_inst|write_reg~q ),
	.datac(!\alt_cal_inst|read~q ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\Selector29~0_combout ),
	.dataf(!\master_write_data[15]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[15]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[15]~7 .extended_lut = "off";
defparam \master_write_data[15]~7 .lut_mask = 64'hD5C0000000000000;
defparam \master_write_data[15]~7 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[15]~8 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.000000~q ),
	.datac(!\Selector1~3_combout ),
	.datad(!\state.ADDRESS_OFFSET_STATE~q ),
	.datae(!\state.WAIT_FOR_NEXT_STATE~q ),
	.dataf(!\Selector45~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[15]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[15]~8 .extended_lut = "off";
defparam \master_write_data[15]~8 .lut_mask = 64'h0000000003000200;
defparam \master_write_data[15]~8 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[15]~9 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.WRITE_DATA_STATE~q ),
	.datae(!\master_write_data[7]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[15]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[15]~9 .extended_lut = "off";
defparam \master_write_data[15]~9 .lut_mask = 64'h0000FF040000FF04;
defparam \master_write_data[15]~9 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[15]~10 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!\state.CHECK_PMUTEX_STATE~q ),
	.datac(!\master_write_data[15]~5_combout ),
	.datad(!\master_write_data[15]~7_combout ),
	.datae(!\master_write_data[15]~8_combout ),
	.dataf(!\master_write_data[15]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[15]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[15]~10 .extended_lut = "off";
defparam \master_write_data[15]~10 .lut_mask = 64'h00000000DD1DFFFF;
defparam \master_write_data[15]~10 .shared_arith = "off";

cyclonev_lcell_comb \Selector67~2 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.GET_TESTBUS_ADDR_STATE~q ),
	.datac(!\Selector77~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector67~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector67~2 .extended_lut = "off";
defparam \Selector67~2 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \Selector67~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector67~1 (
	.dataa(!\master_write~0_combout ),
	.datab(!\state.WRITE_DATA_STATE~q ),
	.datac(!\alt_cal_inst|dataout[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector67~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector67~1 .extended_lut = "off";
defparam \Selector67~1 .lut_mask = 64'h0101010101010101;
defparam \Selector67~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector67~3 (
	.dataa(!\Selector38~0_combout ),
	.datab(!\Selector67~2_combout ),
	.datac(!\Selector67~0_combout ),
	.datad(!\Selector67~1_combout ),
	.datae(!\Selector46~1_combout ),
	.dataf(!master_write_data_11),
	.datag(!\master_write~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector67~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector67~3 .extended_lut = "on";
defparam \Selector67~3 .lut_mask = 64'h5FFF55FFFFFFF7FF;
defparam \Selector67~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector66~0 (
	.dataa(!\state.WRITE_DATA_STATE~q ),
	.datab(!\state.ADDRESS_OFFSET_STATE~q ),
	.datac(!\alt_cal_inst|alt_cal_channel[0]~q ),
	.datad(!\alt_cal_inst|dataout[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector66~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector66~0 .extended_lut = "off";
defparam \Selector66~0 .lut_mask = 64'h0257025702570257;
defparam \Selector66~0 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[12]~11 (
	.dataa(!\alt_cal_inst|alt_cal_busy~q ),
	.datab(!\state.000000~q ),
	.datac(!\Selector1~3_combout ),
	.datad(!\state.WAIT_FOR_NEXT_STATE~q ),
	.datae(!\Selector45~8_combout ),
	.dataf(!\Selector38~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[12]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[12]~11 .extended_lut = "off";
defparam \master_write_data[12]~11 .lut_mask = 64'hFFFFFCFD00000000;
defparam \master_write_data[12]~11 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[12]~12 (
	.dataa(!mutex_grant),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.WRITE_DATA_STATE~q ),
	.datae(!\state.ADDRESS_OFFSET_STATE~q ),
	.dataf(!\master_write_data[7]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[12]~12 .extended_lut = "off";
defparam \master_write_data[12]~12 .lut_mask = 64'h00000000FF040404;
defparam \master_write_data[12]~12 .shared_arith = "off";

cyclonev_lcell_comb \master_write_data[12]~13 (
	.dataa(!\master_write~0_combout ),
	.datab(!\Selector1~3_combout ),
	.datac(!\state.CHECK_PMUTEX_STATE~q ),
	.datad(!\master_write_data[15]~7_combout ),
	.datae(!\master_write_data[12]~11_combout ),
	.dataf(!\master_write_data[12]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_write_data[12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_write_data[12]~13 .extended_lut = "off";
defparam \master_write_data[12]~13 .lut_mask = 64'h00000000FFFFF040;
defparam \master_write_data[12]~13 .shared_arith = "off";

cyclonev_lcell_comb \Selector65~0 (
	.dataa(!\state.WRITE_DATA_STATE~q ),
	.datab(!\state.ADDRESS_OFFSET_STATE~q ),
	.datac(!\alt_cal_inst|alt_cal_channel[1]~q ),
	.datad(!\alt_cal_inst|dataout[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector65~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector65~0 .extended_lut = "off";
defparam \Selector65~0 .lut_mask = 64'h0257025702570257;
defparam \Selector65~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector64~0 (
	.dataa(!\state.WRITE_DATA_STATE~q ),
	.datab(!\alt_cal_inst|dataout[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector64~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector64~0 .extended_lut = "off";
defparam \Selector64~0 .lut_mask = 64'h1111111111111111;
defparam \Selector64~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector63~0 (
	.dataa(!\state.WRITE_DATA_STATE~q ),
	.datab(!\alt_cal_inst|dataout[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector63~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector63~0 .extended_lut = "off";
defparam \Selector63~0 .lut_mask = 64'h1111111111111111;
defparam \Selector63~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_arbiter_acq_3 (
	grant_0,
	req_and_use_mutex,
	mutex_grant)/* synthesis synthesis_greybox=0 */;
input 	grant_0;
input 	req_and_use_mutex;
output 	mutex_grant;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \mutex_grant~0 (
	.dataa(!grant_0),
	.datab(!req_and_use_mutex),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mutex_grant),
	.sumout(),
	.cout(),
	.shareout());
defparam \mutex_grant~0 .extended_lut = "off";
defparam \mutex_grant~0 .lut_mask = 64'h1111111111111111;
defparam \mutex_grant~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_cal_av_1 (
	alt_cal_busy1,
	write_reg1,
	read1,
	alt_cal_channel_9,
	alt_cal_channel_6,
	alt_cal_channel_7,
	alt_cal_channel_8,
	alt_cal_channel_0,
	alt_cal_channel_1,
	alt_cal_channel_2,
	alt_cal_channel_3,
	alt_cal_channel_4,
	alt_cal_channel_5,
	alt_cal_remap_addr_2,
	alt_cal_remap_addr_7,
	alt_cal_remap_addr_10,
	alt_cal_remap_addr_8,
	alt_cal_remap_addr_9,
	alt_cal_remap_addr_1,
	alt_cal_remap_addr_0,
	alt_cal_remap_addr_11,
	alt_cal_remap_addr_3,
	alt_cal_remap_addr_4,
	alt_cal_remap_addr_5,
	alt_cal_remap_addr_6,
	address_1,
	address_0,
	address_4,
	reset,
	start,
	start0q,
	alt_cal_dprio_busy,
	dataout_1,
	dataout_2,
	dataout_0,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_15,
	alt_cal_dprio_datain_14,
	alt_cal_dprio_datain_1,
	alt_cal_dprio_datain_0,
	alt_cal_dprio_datain_3,
	alt_cal_dprio_datain_4,
	alt_cal_dprio_datain_5,
	alt_cal_dprio_datain_6,
	alt_cal_dprio_datain_7,
	alt_cal_dprio_datain_8,
	alt_cal_dprio_datain_9,
	alt_cal_dprio_datain_10,
	alt_cal_dprio_datain_11,
	alt_cal_dprio_datain_12,
	alt_cal_dprio_datain_13,
	alt_cal_dprio_datain_15,
	out_narrow_0,
	out_narrow_1,
	out_narrow_2,
	out_narrow_3,
	clock)/* synthesis synthesis_greybox=0 */;
output 	alt_cal_busy1;
output 	write_reg1;
output 	read1;
output 	alt_cal_channel_9;
output 	alt_cal_channel_6;
output 	alt_cal_channel_7;
output 	alt_cal_channel_8;
output 	alt_cal_channel_0;
output 	alt_cal_channel_1;
output 	alt_cal_channel_2;
output 	alt_cal_channel_3;
output 	alt_cal_channel_4;
output 	alt_cal_channel_5;
input 	alt_cal_remap_addr_2;
input 	alt_cal_remap_addr_7;
input 	alt_cal_remap_addr_10;
input 	alt_cal_remap_addr_8;
input 	alt_cal_remap_addr_9;
input 	alt_cal_remap_addr_1;
input 	alt_cal_remap_addr_0;
input 	alt_cal_remap_addr_11;
input 	alt_cal_remap_addr_3;
input 	alt_cal_remap_addr_4;
input 	alt_cal_remap_addr_5;
input 	alt_cal_remap_addr_6;
output 	address_1;
output 	address_0;
output 	address_4;
input 	reset;
input 	start;
input 	start0q;
input 	alt_cal_dprio_busy;
output 	dataout_1;
output 	dataout_2;
output 	dataout_0;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_15;
input 	alt_cal_dprio_datain_14;
input 	alt_cal_dprio_datain_1;
input 	alt_cal_dprio_datain_0;
input 	alt_cal_dprio_datain_3;
input 	alt_cal_dprio_datain_4;
input 	alt_cal_dprio_datain_5;
input 	alt_cal_dprio_datain_6;
input 	alt_cal_dprio_datain_7;
input 	alt_cal_dprio_datain_8;
input 	alt_cal_dprio_datain_9;
input 	alt_cal_dprio_datain_10;
input 	alt_cal_dprio_datain_11;
input 	alt_cal_dprio_datain_12;
input 	alt_cal_dprio_datain_13;
input 	alt_cal_dprio_datain_15;
input 	out_narrow_0;
input 	out_narrow_1;
input 	out_narrow_2;
input 	out_narrow_3;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pd0_det|ff2~q ;
wire \pd90_det|ff2~q ;
wire \pd180_det|ff2~q ;
wire \pd270_det|ff2~q ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \LessThan1~2_combout ;
wire \Equal11~0_combout ;
wire \Equal11~1_combout ;
wire \Equal11~2_combout ;
wire \Selector74~0_combout ;
wire \done~q ;
wire \p0addr~q ;
wire \Selector11~0_combout ;
wire \Selector12~0_combout ;
wire \Selector12~1_combout ;
wire \state.CH_WAIT~q ;
wire \Add4~5_sumout ;
wire \Add4~2 ;
wire \Add4~17_sumout ;
wire \Equal1~0_combout ;
wire \Selector56~0_combout ;
wire \ch_testbus0q[0]~q ;
wire \ch_testbus1q[0]~q ;
wire \pd_0~0_combout ;
wire \Equal0~1_combout ;
wire \Selector86~0_combout ;
wire \ret_state.PDOF_TEST_RD~q ;
wire \Selector20~0_combout ;
wire \state.PDOF_TEST_RD~q ;
wire \Selector81~0_combout ;
wire \Selector82~0_combout ;
wire \Selector84~0_combout ;
wire \ret_state.DPRIO_WAIT~q ;
wire \Selector15~0_combout ;
wire \state.DPRIO_WAIT~q ;
wire \pd_0[0]~1_combout ;
wire \pd_0[0]~q ;
wire \pd_0_p[0]~1_combout ;
wire \pd_0_p[0]~q ;
wire \pd_1~0_combout ;
wire \pd_1[0]~q ;
wire \pd_1_p[0]~q ;
wire \WideOr8~0_combout ;
wire \recal_counter[0]~0_combout ;
wire \recal_counter[0]~1_combout ;
wire \recal_counter[0]~q ;
wire \Add5~0_combout ;
wire \recal_counter[1]~q ;
wire \Selector57~2_combout ;
wire \cal_pd0_l~0_combout ;
wire \Selector56~3_combout ;
wire \cal_pd0_l[0]~1_combout ;
wire \cal_pd0_l[3]~q ;
wire \cal_pd0_l~4_combout ;
wire \cal_pd0_l[2]~q ;
wire \cal_pd0_l~3_combout ;
wire \cal_pd0_l[1]~q ;
wire \cal_pd0_l~2_combout ;
wire \cal_pd0_l[0]~q ;
wire \Add0~18_cout ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \cal_pd0~0_combout ;
wire \cal_pd0~3_combout ;
wire \cal_pd0~6_combout ;
wire \Selector24~0_combout ;
wire \cal_pd0[1]~q ;
wire \Add6~1_combout ;
wire \Add0~6 ;
wire \Add0~13_sumout ;
wire \cal_pd0~5_combout ;
wire \Selector23~0_combout ;
wire \cal_pd0[2]~q ;
wire \Equal4~0_combout ;
wire \Selector65~0_combout ;
wire \Selector65~1_combout ;
wire \ignore_solid[0]~q ;
wire \data_e0q[0]~q ;
wire \data_e1q[0]~q ;
wire \cal_pd0~1_combout ;
wire \Selector61~0_combout ;
wire \cal_inc[0]~q ;
wire \cal_pd0~2_combout ;
wire \Add0~9_sumout ;
wire \Selector25~0_combout ;
wire \Selector25~1_combout ;
wire \Selector25~2_combout ;
wire \cal_pd0[0]~q ;
wire \Add6~0_combout ;
wire \Add0~14 ;
wire \Add0~1_sumout ;
wire \cal_pd0~4_combout ;
wire \Selector22~0_combout ;
wire \cal_pd0[3]~q ;
wire \Selector57~0_combout ;
wire \Selector57~1_combout ;
wire \cal_done[0]~q ;
wire \ch_testbus0q[1]~q ;
wire \ch_testbus1q[1]~q ;
wire \pd_0~2_combout ;
wire \pd_0[1]~q ;
wire \pd_0_p[1]~q ;
wire \pd_1~1_combout ;
wire \pd_1[1]~q ;
wire \pd_1_p[1]~q ;
wire \cal_pd90_l~0_combout ;
wire \cal_pd90_l[3]~1_combout ;
wire \cal_pd90_l[3]~q ;
wire \cal_pd90~2_combout ;
wire \cal_pd90~0_combout ;
wire \cal_pd90_l~3_combout ;
wire \cal_pd90_l[1]~q ;
wire \cal_pd90_l~2_combout ;
wire \cal_pd90_l[0]~q ;
wire \Add1~18_cout ;
wire \Add1~5_sumout ;
wire \Selector29~0_combout ;
wire \Selector29~1_combout ;
wire \Selector29~2_combout ;
wire \cal_pd90[0]~q ;
wire \cal_pd90_l~4_combout ;
wire \cal_pd90_l[2]~q ;
wire \Equal6~0_combout ;
wire \Selector64~0_combout ;
wire \Selector64~1_combout ;
wire \ignore_solid[1]~q ;
wire \data_e0q[1]~q ;
wire \data_e1q[1]~q ;
wire \cal_pd90~1_combout ;
wire \Selector60~0_combout ;
wire \cal_inc[1]~q ;
wire \Add1~6 ;
wire \Add1~13_sumout ;
wire \cal_pd90~3_combout ;
wire \cal_pd90~6_combout ;
wire \Selector28~0_combout ;
wire \cal_pd90[1]~q ;
wire \Add7~1_combout ;
wire \Add1~14 ;
wire \Add1~9_sumout ;
wire \cal_pd90~5_combout ;
wire \Selector27~0_combout ;
wire \cal_pd90[2]~q ;
wire \Add7~0_combout ;
wire \Add1~10 ;
wire \Add1~1_sumout ;
wire \cal_pd90~4_combout ;
wire \Selector26~0_combout ;
wire \cal_pd90[3]~q ;
wire \Selector56~1_combout ;
wire \Selector56~2_combout ;
wire \cal_done[1]~q ;
wire \ch_testbus0q[2]~q ;
wire \ch_testbus1q[2]~q ;
wire \pd_0~3_combout ;
wire \pd_0[2]~q ;
wire \pd_0_p[2]~q ;
wire \pd_1~2_combout ;
wire \pd_1[2]~q ;
wire \pd_1_p[2]~q ;
wire \cal_pd180_l~0_combout ;
wire \cal_pd180_l[3]~1_combout ;
wire \cal_pd180_l[3]~q ;
wire \cal_pd180~2_combout ;
wire \cal_pd180~0_combout ;
wire \cal_pd180_l~3_combout ;
wire \cal_pd180_l[1]~q ;
wire \cal_pd180_l~2_combout ;
wire \cal_pd180_l[0]~q ;
wire \Add2~18_cout ;
wire \Add2~5_sumout ;
wire \Selector33~0_combout ;
wire \Selector33~1_combout ;
wire \Selector33~2_combout ;
wire \cal_pd180[0]~q ;
wire \cal_pd180_l~4_combout ;
wire \cal_pd180_l[2]~q ;
wire \Equal8~0_combout ;
wire \Selector63~0_combout ;
wire \Selector63~1_combout ;
wire \ignore_solid[2]~q ;
wire \data_e0q[2]~q ;
wire \data_e1q[2]~q ;
wire \cal_pd180~1_combout ;
wire \Selector59~0_combout ;
wire \cal_inc[2]~q ;
wire \Add2~6 ;
wire \Add2~13_sumout ;
wire \cal_pd180~3_combout ;
wire \cal_pd180~6_combout ;
wire \Selector32~0_combout ;
wire \cal_pd180[1]~q ;
wire \Add8~1_combout ;
wire \Add2~14 ;
wire \Add2~9_sumout ;
wire \cal_pd180~5_combout ;
wire \Selector31~0_combout ;
wire \cal_pd180[2]~q ;
wire \Add8~0_combout ;
wire \Add2~10 ;
wire \Add2~1_sumout ;
wire \cal_pd180~4_combout ;
wire \Selector30~0_combout ;
wire \cal_pd180[3]~q ;
wire \Selector55~0_combout ;
wire \Selector55~1_combout ;
wire \cal_done[2]~q ;
wire \ch_testbus0q[3]~q ;
wire \ch_testbus1q[3]~q ;
wire \pd_0~4_combout ;
wire \pd_0[3]~q ;
wire \pd_0_p[3]~q ;
wire \pd_1~3_combout ;
wire \pd_1[3]~q ;
wire \pd_1_p[3]~q ;
wire \Selector58~0_combout ;
wire \cal_inc[3]~q ;
wire \cal_pd270_l~0_combout ;
wire \cal_pd270_l[1]~1_combout ;
wire \cal_pd270_l[3]~q ;
wire \Add9~1_combout ;
wire \cal_pd270_l~4_combout ;
wire \cal_pd270_l[2]~q ;
wire \cal_pd270_l~3_combout ;
wire \cal_pd270_l[1]~q ;
wire \cal_pd270_l~2_combout ;
wire \cal_pd270_l[0]~q ;
wire \Add3~18_cout ;
wire \Add3~2 ;
wire \Add3~14 ;
wire \Add3~9_sumout ;
wire \Selector35~0_combout ;
wire \Selector35~1_combout ;
wire \cal_pd270[2]~q ;
wire \cal_pd270~1_combout ;
wire \cal_pd270~2_combout ;
wire \Add9~2_combout ;
wire \Add3~13_sumout ;
wire \Selector36~0_combout ;
wire \Selector36~1_combout ;
wire \cal_pd270[1]~q ;
wire \Add3~1_sumout ;
wire \Selector37~0_combout ;
wire \cal_pd270[0]~q ;
wire \Equal10~0_combout ;
wire \cal_pd270~0_combout ;
wire \Add9~0_combout ;
wire \Add3~10 ;
wire \Add3~5_sumout ;
wire \Selector34~0_combout ;
wire \Selector34~1_combout ;
wire \cal_pd270[3]~q ;
wire \Selector62~0_combout ;
wire \Selector62~1_combout ;
wire \ignore_solid[3]~q ;
wire \data_e0q[3]~q ;
wire \data_e1q[3]~q ;
wire \edges[3]~0_combout ;
wire \Selector54~0_combout ;
wire \cal_done[3]~q ;
wire \WideAnd0~combout ;
wire \Selector0~0_combout ;
wire \cal_en~q ;
wire \Selector83~0_combout ;
wire \ret_state.CAL_PD_WR~q ;
wire \Selector14~0_combout ;
wire \state.CAL_PD_WR~q ;
wire \WideAnd1~0_combout ;
wire \WideAnd1~1_combout ;
wire \WideAnd2~0_combout ;
wire \WideAnd3~0_combout ;
wire \WideAnd4~0_combout ;
wire \Selector75~0_combout ;
wire \Selector75~1_combout ;
wire \Selector75~2_combout ;
wire \Selector75~3_combout ;
wire \do_recal~q ;
wire \always1~0_combout ;
wire \counter[2]~1_combout ;
wire \counter[3]~q ;
wire \Add4~18 ;
wire \Add4~13_sumout ;
wire \counter[4]~q ;
wire \Add4~14 ;
wire \Add4~29_sumout ;
wire \counter[5]~q ;
wire \Add4~30 ;
wire \Add4~25_sumout ;
wire \counter[6]~q ;
wire \pd_0_p[0]~0_combout ;
wire \counter[2]~0_combout ;
wire \counter[0]~q ;
wire \Add4~6 ;
wire \Add4~21_sumout ;
wire \counter[1]~q ;
wire \Add4~22 ;
wire \Add4~1_sumout ;
wire \counter[2]~q ;
wire \Add4~26 ;
wire \Add4~9_sumout ;
wire \counter[7]~q ;
wire \Equal0~0_combout ;
wire \Equal1~1_combout ;
wire \Selector16~0_combout ;
wire \state.SAMPLE_TB~q ;
wire \state~30_combout ;
wire \state.TEST_INPUT~q ;
wire \Selector13~0_combout ;
wire \state.TESTBUS_SET~q ;
wire \state~29_combout ;
wire \state.CHECK_PLL_RD~q ;
wire \Selector18~0_combout ;
wire \Selector18~1_combout ;
wire \state.DPRIO_READ~q ;
wire \state~25_combout ;
wire \Selector87~0_combout ;
wire \ret_state.PDOF_TEST_WR~q ;
wire \Selector21~0_combout ;
wire \state.PDOF_TEST_WR~q ;
wire \Selector104~0_combout ;
wire \Selector19~0_combout ;
wire \state.DPRIO_WRITE~q ;
wire \Selector82~1_combout ;
wire \did_dprio~q ;
wire \state~28_combout ;
wire \Selector17~0_combout ;
wire \Selector17~1_combout ;
wire \Selector85~0_combout ;
wire \ret_state.CH_ADV~q ;
wire \Selector17~2_combout ;
wire \Selector17~3_combout ;
wire \state.CH_ADV~q ;
wire \ret_state~12_combout ;
wire \ret_state.IDLE~q ;
wire \state~26_combout ;
wire \state~27_combout ;
wire \state.IDLE~q ;
wire \alt_cal_busy~0_combout ;
wire \Selector104~1_combout ;
wire \Selector81~1_combout ;
wire \Add10~18 ;
wire \Add10~22 ;
wire \Add10~26 ;
wire \Add10~30 ;
wire \Add10~34 ;
wire \Add10~38 ;
wire \Add10~6 ;
wire \Add10~10 ;
wire \Add10~14 ;
wire \Add10~1_sumout ;
wire \Selector1~0_combout ;
wire \Selector10~0_combout ;
wire \Add10~5_sumout ;
wire \Selector4~0_combout ;
wire \Add10~9_sumout ;
wire \Selector3~0_combout ;
wire \Add10~13_sumout ;
wire \Selector2~0_combout ;
wire \Add10~17_sumout ;
wire \Selector10~1_combout ;
wire \Add10~21_sumout ;
wire \Selector9~0_combout ;
wire \Add10~25_sumout ;
wire \Selector8~0_combout ;
wire \Add10~29_sumout ;
wire \Selector7~0_combout ;
wire \Add10~33_sumout ;
wire \Selector6~0_combout ;
wire \Add10~37_sumout ;
wire \Selector5~0_combout ;
wire \Selector79~0_combout ;
wire \Selector80~0_combout ;
wire \Selector76~0_combout ;
wire \dataout[0]~0_combout ;
wire \dataout~1_combout ;
wire \dataout[0]~2_combout ;
wire \dataout~3_combout ;
wire \dataout~4_combout ;
wire \dataout~5_combout ;
wire \dataout[5]~6_combout ;
wire \dataout~7_combout ;
wire \dataout~8_combout ;
wire \dataout~9_combout ;
wire \dataout~10_combout ;
wire \dataout[8]~11_combout ;
wire \dataout~12_combout ;
wire \dataout~13_combout ;
wire \dataout~14_combout ;
wire \dataout~15_combout ;
wire \dataout[13]~16_combout ;
wire \dataout~17_combout ;
wire \dataout~18_combout ;
wire \dataout~19_combout ;
wire \dataout~20_combout ;


RECONFIGURE_IP_alt_cal_edge_detect_2 pd270_det(
	.reset(\state.DPRIO_WRITE~q ),
	.ff21(\pd270_det|ff2~q ),
	.testbus(out_narrow_3));

RECONFIGURE_IP_alt_cal_edge_detect_1 pd180_det(
	.reset(\state.DPRIO_WRITE~q ),
	.ff21(\pd180_det|ff2~q ),
	.testbus(out_narrow_2));

RECONFIGURE_IP_alt_cal_edge_detect_3 pd90_det(
	.reset(\state.DPRIO_WRITE~q ),
	.ff21(\pd90_det|ff2~q ),
	.testbus(out_narrow_1));

RECONFIGURE_IP_alt_cal_edge_detect pd0_det(
	.reset(\state.DPRIO_WRITE~q ),
	.ff21(\pd0_det|ff2~q ),
	.testbus(out_narrow_0));

dffeas alt_cal_busy(
	.clk(clock),
	.d(\alt_cal_busy~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_busy1),
	.prn(vcc));
defparam alt_cal_busy.is_wysiwyg = "true";
defparam alt_cal_busy.power_up = "low";

dffeas write_reg(
	.clk(clock),
	.d(\Selector104~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(write_reg1),
	.prn(vcc));
defparam write_reg.is_wysiwyg = "true";
defparam write_reg.power_up = "low";

dffeas read(
	.clk(clock),
	.d(\Selector81~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(read1),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas \alt_cal_channel[9] (
	.clk(clock),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_9),
	.prn(vcc));
defparam \alt_cal_channel[9] .is_wysiwyg = "true";
defparam \alt_cal_channel[9] .power_up = "low";

dffeas \alt_cal_channel[6] (
	.clk(clock),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_6),
	.prn(vcc));
defparam \alt_cal_channel[6] .is_wysiwyg = "true";
defparam \alt_cal_channel[6] .power_up = "low";

dffeas \alt_cal_channel[7] (
	.clk(clock),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_7),
	.prn(vcc));
defparam \alt_cal_channel[7] .is_wysiwyg = "true";
defparam \alt_cal_channel[7] .power_up = "low";

dffeas \alt_cal_channel[8] (
	.clk(clock),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_8),
	.prn(vcc));
defparam \alt_cal_channel[8] .is_wysiwyg = "true";
defparam \alt_cal_channel[8] .power_up = "low";

dffeas \alt_cal_channel[0] (
	.clk(clock),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_0),
	.prn(vcc));
defparam \alt_cal_channel[0] .is_wysiwyg = "true";
defparam \alt_cal_channel[0] .power_up = "low";

dffeas \alt_cal_channel[1] (
	.clk(clock),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_1),
	.prn(vcc));
defparam \alt_cal_channel[1] .is_wysiwyg = "true";
defparam \alt_cal_channel[1] .power_up = "low";

dffeas \alt_cal_channel[2] (
	.clk(clock),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_2),
	.prn(vcc));
defparam \alt_cal_channel[2] .is_wysiwyg = "true";
defparam \alt_cal_channel[2] .power_up = "low";

dffeas \alt_cal_channel[3] (
	.clk(clock),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_3),
	.prn(vcc));
defparam \alt_cal_channel[3] .is_wysiwyg = "true";
defparam \alt_cal_channel[3] .power_up = "low";

dffeas \alt_cal_channel[4] (
	.clk(clock),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_4),
	.prn(vcc));
defparam \alt_cal_channel[4] .is_wysiwyg = "true";
defparam \alt_cal_channel[4] .power_up = "low";

dffeas \alt_cal_channel[5] (
	.clk(clock),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(alt_cal_channel_5),
	.prn(vcc));
defparam \alt_cal_channel[5] .is_wysiwyg = "true";
defparam \alt_cal_channel[5] .power_up = "low";

dffeas \address[1] (
	.clk(clock),
	.d(\Selector79~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(address_1),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[0] (
	.clk(clock),
	.d(\Selector80~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(address_0),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[4] (
	.clk(clock),
	.d(\Selector76~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(address_4),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \dataout[1] (
	.clk(clock),
	.d(\dataout~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_1),
	.prn(vcc));
defparam \dataout[1] .is_wysiwyg = "true";
defparam \dataout[1] .power_up = "low";

dffeas \dataout[2] (
	.clk(clock),
	.d(\dataout~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_2),
	.prn(vcc));
defparam \dataout[2] .is_wysiwyg = "true";
defparam \dataout[2] .power_up = "low";

dffeas \dataout[0] (
	.clk(clock),
	.d(\dataout~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_0),
	.prn(vcc));
defparam \dataout[0] .is_wysiwyg = "true";
defparam \dataout[0] .power_up = "low";

dffeas \dataout[3] (
	.clk(clock),
	.d(\dataout~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_3),
	.prn(vcc));
defparam \dataout[3] .is_wysiwyg = "true";
defparam \dataout[3] .power_up = "low";

dffeas \dataout[4] (
	.clk(clock),
	.d(\dataout~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_4),
	.prn(vcc));
defparam \dataout[4] .is_wysiwyg = "true";
defparam \dataout[4] .power_up = "low";

dffeas \dataout[5] (
	.clk(clock),
	.d(\dataout~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_5),
	.prn(vcc));
defparam \dataout[5] .is_wysiwyg = "true";
defparam \dataout[5] .power_up = "low";

dffeas \dataout[6] (
	.clk(clock),
	.d(\dataout~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_6),
	.prn(vcc));
defparam \dataout[6] .is_wysiwyg = "true";
defparam \dataout[6] .power_up = "low";

dffeas \dataout[7] (
	.clk(clock),
	.d(\dataout~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_7),
	.prn(vcc));
defparam \dataout[7] .is_wysiwyg = "true";
defparam \dataout[7] .power_up = "low";

dffeas \dataout[8] (
	.clk(clock),
	.d(\dataout~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_8),
	.prn(vcc));
defparam \dataout[8] .is_wysiwyg = "true";
defparam \dataout[8] .power_up = "low";

dffeas \dataout[9] (
	.clk(clock),
	.d(\dataout~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_9),
	.prn(vcc));
defparam \dataout[9] .is_wysiwyg = "true";
defparam \dataout[9] .power_up = "low";

dffeas \dataout[10] (
	.clk(clock),
	.d(\dataout~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_10),
	.prn(vcc));
defparam \dataout[10] .is_wysiwyg = "true";
defparam \dataout[10] .power_up = "low";

dffeas \dataout[11] (
	.clk(clock),
	.d(\dataout~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_11),
	.prn(vcc));
defparam \dataout[11] .is_wysiwyg = "true";
defparam \dataout[11] .power_up = "low";

dffeas \dataout[12] (
	.clk(clock),
	.d(\dataout~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_12),
	.prn(vcc));
defparam \dataout[12] .is_wysiwyg = "true";
defparam \dataout[12] .power_up = "low";

dffeas \dataout[13] (
	.clk(clock),
	.d(\dataout~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_13),
	.prn(vcc));
defparam \dataout[13] .is_wysiwyg = "true";
defparam \dataout[13] .power_up = "low";

dffeas \dataout[14] (
	.clk(clock),
	.d(\dataout~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_14),
	.prn(vcc));
defparam \dataout[14] .is_wysiwyg = "true";
defparam \dataout[14] .power_up = "low";

dffeas \dataout[15] (
	.clk(clock),
	.d(\dataout~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dataout[0]~2_combout ),
	.q(dataout_15),
	.prn(vcc));
defparam \dataout[15] .is_wysiwyg = "true";
defparam \dataout[15] .power_up = "low";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!alt_cal_channel_0),
	.datab(!alt_cal_channel_1),
	.datac(!alt_cal_channel_5),
	.datad(!alt_cal_channel_7),
	.datae(!alt_cal_channel_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h8000000080000000;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!alt_cal_channel_2),
	.datab(!alt_cal_channel_3),
	.datac(!alt_cal_channel_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'h8080808080808080;
defparam \LessThan1~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~2 (
	.dataa(!alt_cal_channel_6),
	.datab(!\LessThan1~0_combout ),
	.datac(!\LessThan1~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~2 .extended_lut = "off";
defparam \LessThan1~2 .lut_mask = 64'h0202020202020202;
defparam \LessThan1~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal11~0 (
	.dataa(!alt_cal_remap_addr_8),
	.datab(!alt_cal_remap_addr_9),
	.datac(!alt_cal_remap_addr_1),
	.datad(!alt_cal_remap_addr_0),
	.datae(!alt_cal_remap_addr_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal11~0 .extended_lut = "off";
defparam \Equal11~0 .lut_mask = 64'h0000000100000001;
defparam \Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal11~1 (
	.dataa(!alt_cal_remap_addr_3),
	.datab(!alt_cal_remap_addr_4),
	.datac(!alt_cal_remap_addr_5),
	.datad(!alt_cal_remap_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal11~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal11~1 .extended_lut = "off";
defparam \Equal11~1 .lut_mask = 64'h0001000100010001;
defparam \Equal11~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal11~2 (
	.dataa(!alt_cal_remap_addr_2),
	.datab(!alt_cal_remap_addr_7),
	.datac(!alt_cal_remap_addr_10),
	.datad(!\Equal11~0_combout ),
	.datae(!\Equal11~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal11~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal11~2 .extended_lut = "off";
defparam \Equal11~2 .lut_mask = 64'h0000000100000001;
defparam \Equal11~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector74~0 (
	.dataa(!alt_cal_channel_9),
	.datab(!\done~q ),
	.datac(!\LessThan1~2_combout ),
	.datad(!\state.CH_ADV~q ),
	.datae(!\state.CH_WAIT~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector74~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector74~0 .extended_lut = "off";
defparam \Selector74~0 .lut_mask = 64'h33F700F733F700F7;
defparam \Selector74~0 .shared_arith = "off";

dffeas done(
	.clk(clock),
	.d(\Selector74~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\done~q ),
	.prn(vcc));
defparam done.is_wysiwyg = "true";
defparam done.power_up = "low";

dffeas p0addr(
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\p0addr~q ),
	.prn(vcc));
defparam p0addr.is_wysiwyg = "true";
defparam p0addr.power_up = "low";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!start),
	.datab(!start0q),
	.datac(!\done~q ),
	.datad(!\p0addr~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h44F444F444F444F4;
defparam \Selector11~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!alt_cal_channel_6),
	.datab(!alt_cal_channel_9),
	.datac(!\LessThan1~0_combout ),
	.datad(!\LessThan1~1_combout ),
	.datae(!\state.CH_ADV~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'h0000000800000008;
defparam \Selector12~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~1 (
	.dataa(!\state.IDLE~q ),
	.datab(!\Selector11~0_combout ),
	.datac(!\Selector12~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~1 .extended_lut = "off";
defparam \Selector12~1 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \Selector12~1 .shared_arith = "off";

dffeas \state.CH_WAIT (
	.clk(clock),
	.d(\Selector12~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CH_WAIT~q ),
	.prn(vcc));
defparam \state.CH_WAIT .is_wysiwyg = "true";
defparam \state.CH_WAIT .power_up = "low";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!\counter[1]~q ),
	.datab(!\counter[6]~q ),
	.datac(!\counter[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0202020202020202;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector56~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\state.SAMPLE_TB~q ),
	.datad(!\always1~0_combout ),
	.datae(!\Equal0~0_combout ),
	.dataf(!\Equal1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector56~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector56~0 .extended_lut = "off";
defparam \Selector56~0 .lut_mask = 64'h404040404040404C;
defparam \Selector56~0 .shared_arith = "off";

dffeas \ch_testbus0q[0] (
	.clk(clock),
	.d(out_narrow_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus0q[0]~q ),
	.prn(vcc));
defparam \ch_testbus0q[0] .is_wysiwyg = "true";
defparam \ch_testbus0q[0] .power_up = "low";

dffeas \ch_testbus1q[0] (
	.clk(clock),
	.d(\ch_testbus0q[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus1q[0]~q ),
	.prn(vcc));
defparam \ch_testbus1q[0] .is_wysiwyg = "true";
defparam \ch_testbus1q[0] .power_up = "low";

cyclonev_lcell_comb \pd_0~0 (
	.dataa(!\pd_0[0]~q ),
	.datab(!\ch_testbus1q[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_0~0 .extended_lut = "off";
defparam \pd_0~0 .lut_mask = 64'h4444444444444444;
defparam \pd_0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\counter[1]~q ),
	.datab(!\counter[6]~q ),
	.datac(!\counter[5]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h0040004000400040;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector86~0 (
	.dataa(!\state.CHECK_PLL_RD~q ),
	.datab(!\Selector82~0_combout ),
	.datac(!\ret_state.PDOF_TEST_RD~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector86~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector86~0 .extended_lut = "off";
defparam \Selector86~0 .lut_mask = 64'h5757575757575757;
defparam \Selector86~0 .shared_arith = "off";

dffeas \ret_state.PDOF_TEST_RD (
	.clk(clock),
	.d(\Selector86~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ret_state.PDOF_TEST_RD~q ),
	.prn(vcc));
defparam \ret_state.PDOF_TEST_RD .is_wysiwyg = "true";
defparam \ret_state.PDOF_TEST_RD .power_up = "low";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!\state~25_combout ),
	.datab(!\ret_state.PDOF_TEST_RD~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h1111111111111111;
defparam \Selector20~0 .shared_arith = "off";

dffeas \state.PDOF_TEST_RD (
	.clk(clock),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.PDOF_TEST_RD~q ),
	.prn(vcc));
defparam \state.PDOF_TEST_RD .is_wysiwyg = "true";
defparam \state.PDOF_TEST_RD .power_up = "low";

cyclonev_lcell_comb \Selector81~0 (
	.dataa(!\state.CHECK_PLL_RD~q ),
	.datab(!\state.PDOF_TEST_RD~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector81~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector81~0 .extended_lut = "off";
defparam \Selector81~0 .lut_mask = 64'h8888888888888888;
defparam \Selector81~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector82~0 (
	.dataa(!\Selector104~0_combout ),
	.datab(!\Selector81~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector82~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector82~0 .extended_lut = "off";
defparam \Selector82~0 .lut_mask = 64'h1111111111111111;
defparam \Selector82~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector84~0 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\Selector82~0_combout ),
	.datac(!\ret_state.DPRIO_WAIT~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector84~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector84~0 .extended_lut = "off";
defparam \Selector84~0 .lut_mask = 64'h5757575757575757;
defparam \Selector84~0 .shared_arith = "off";

dffeas \ret_state.DPRIO_WAIT (
	.clk(clock),
	.d(\Selector84~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ret_state.DPRIO_WAIT~q ),
	.prn(vcc));
defparam \ret_state.DPRIO_WAIT .is_wysiwyg = "true";
defparam \ret_state.DPRIO_WAIT .power_up = "low";

cyclonev_lcell_comb \Selector15~0 (
	.dataa(!\state~25_combout ),
	.datab(!\state.DPRIO_WAIT~q ),
	.datac(!\Equal0~1_combout ),
	.datad(!\ret_state.DPRIO_WAIT~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "off";
defparam \Selector15~0 .lut_mask = 64'h3075307530753075;
defparam \Selector15~0 .shared_arith = "off";

dffeas \state.DPRIO_WAIT (
	.clk(clock),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.DPRIO_WAIT~q ),
	.prn(vcc));
defparam \state.DPRIO_WAIT .is_wysiwyg = "true";
defparam \state.DPRIO_WAIT .power_up = "low";

cyclonev_lcell_comb \pd_0[0]~1 (
	.dataa(!reset),
	.datab(!\state.SAMPLE_TB~q ),
	.datac(!\state.DPRIO_WAIT~q ),
	.datad(!\Equal0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_0[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_0[0]~1 .extended_lut = "off";
defparam \pd_0[0]~1 .lut_mask = 64'h1015101510151015;
defparam \pd_0[0]~1 .shared_arith = "off";

dffeas \pd_0[0] (
	.clk(clock),
	.d(\pd_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_0[0]~q ),
	.prn(vcc));
defparam \pd_0[0] .is_wysiwyg = "true";
defparam \pd_0[0] .power_up = "low";

cyclonev_lcell_comb \pd_0_p[0]~1 (
	.dataa(!reset),
	.datab(!\counter[1]~q ),
	.datac(!\counter[6]~q ),
	.datad(!\counter[5]~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(!\state.DPRIO_WAIT~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_0_p[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_0_p[0]~1 .extended_lut = "off";
defparam \pd_0_p[0]~1 .lut_mask = 64'h0000000000001000;
defparam \pd_0_p[0]~1 .shared_arith = "off";

dffeas \pd_0_p[0] (
	.clk(clock),
	.d(\pd_0[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_0_p[0]~q ),
	.prn(vcc));
defparam \pd_0_p[0] .is_wysiwyg = "true";
defparam \pd_0_p[0] .power_up = "low";

cyclonev_lcell_comb \pd_1~0 (
	.dataa(!\pd_1[0]~q ),
	.datab(!\ch_testbus1q[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_1~0 .extended_lut = "off";
defparam \pd_1~0 .lut_mask = 64'h1111111111111111;
defparam \pd_1~0 .shared_arith = "off";

dffeas \pd_1[0] (
	.clk(clock),
	.d(\pd_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_1[0]~q ),
	.prn(vcc));
defparam \pd_1[0] .is_wysiwyg = "true";
defparam \pd_1[0] .power_up = "low";

dffeas \pd_1_p[0] (
	.clk(clock),
	.d(\pd_1[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_1_p[0]~q ),
	.prn(vcc));
defparam \pd_1_p[0] .is_wysiwyg = "true";
defparam \pd_1_p[0] .power_up = "low";

cyclonev_lcell_comb \WideOr8~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\state.SAMPLE_TB~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr8~0 .extended_lut = "off";
defparam \WideOr8~0 .lut_mask = 64'h8080808080808080;
defparam \WideOr8~0 .shared_arith = "off";

cyclonev_lcell_comb \recal_counter[0]~0 (
	.dataa(!reset),
	.datab(!\state.SAMPLE_TB~q ),
	.datac(!\always1~0_combout ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\recal_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \recal_counter[0]~0 .extended_lut = "off";
defparam \recal_counter[0]~0 .lut_mask = 64'hAAAAAAABAAAAAAAB;
defparam \recal_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \recal_counter[0]~1 (
	.dataa(!reset),
	.datab(!\recal_counter[0]~q ),
	.datac(!\recal_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\recal_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \recal_counter[0]~1 .extended_lut = "off";
defparam \recal_counter[0]~1 .lut_mask = 64'h3434343434343434;
defparam \recal_counter[0]~1 .shared_arith = "off";

dffeas \recal_counter[0] (
	.clk(clock),
	.d(\recal_counter[0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\recal_counter[0]~q ),
	.prn(vcc));
defparam \recal_counter[0] .is_wysiwyg = "true";
defparam \recal_counter[0] .power_up = "low";

cyclonev_lcell_comb \Add5~0 (
	.dataa(!\recal_counter[0]~q ),
	.datab(!\recal_counter[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~0 .extended_lut = "off";
defparam \Add5~0 .lut_mask = 64'h6666666666666666;
defparam \Add5~0 .shared_arith = "off";

dffeas \recal_counter[1] (
	.clk(clock),
	.d(\Add5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(\recal_counter[0]~0_combout ),
	.q(\recal_counter[1]~q ),
	.prn(vcc));
defparam \recal_counter[1] .is_wysiwyg = "true";
defparam \recal_counter[1] .power_up = "low";

cyclonev_lcell_comb \Selector57~2 (
	.dataa(!\state.SAMPLE_TB~q ),
	.datab(!\do_recal~q ),
	.datac(!\recal_counter[0]~q ),
	.datad(!\recal_counter[1]~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(!\Equal1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector57~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector57~2 .extended_lut = "off";
defparam \Selector57~2 .lut_mask = 64'h5555555555554445;
defparam \Selector57~2 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd0_l~0 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0_l~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0_l~0 .extended_lut = "off";
defparam \cal_pd0_l~0 .lut_mask = 64'h0101010101010101;
defparam \cal_pd0_l~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector56~3 (
	.dataa(!\state.SAMPLE_TB~q ),
	.datab(!\WideOr8~0_combout ),
	.datac(!\always1~0_combout ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector56~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector56~3 .extended_lut = "off";
defparam \Selector56~3 .lut_mask = 64'h8888888C8888888C;
defparam \Selector56~3 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd0_l[0]~1 (
	.dataa(!reset),
	.datab(!\cal_done[0]~q ),
	.datac(!\state.TEST_INPUT~q ),
	.datad(!\Selector56~3_combout ),
	.datae(!\cal_inc[0]~q ),
	.dataf(!\cal_pd0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0_l[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0_l[0]~1 .extended_lut = "off";
defparam \cal_pd0_l[0]~1 .lut_mask = 64'hAAFEAAFAAAFAAAFA;
defparam \cal_pd0_l[0]~1 .shared_arith = "off";

dffeas \cal_pd0_l[3] (
	.clk(clock),
	.d(\cal_pd0_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd0_l[0]~1_combout ),
	.q(\cal_pd0_l[3]~q ),
	.prn(vcc));
defparam \cal_pd0_l[3] .is_wysiwyg = "true";
defparam \cal_pd0_l[3] .power_up = "low";

cyclonev_lcell_comb \cal_pd0_l~4 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0_l~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0_l~4 .extended_lut = "off";
defparam \cal_pd0_l~4 .lut_mask = 64'h0101010101010101;
defparam \cal_pd0_l~4 .shared_arith = "off";

dffeas \cal_pd0_l[2] (
	.clk(clock),
	.d(\cal_pd0_l~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd0_l[0]~1_combout ),
	.q(\cal_pd0_l[2]~q ),
	.prn(vcc));
defparam \cal_pd0_l[2] .is_wysiwyg = "true";
defparam \cal_pd0_l[2] .power_up = "low";

cyclonev_lcell_comb \cal_pd0_l~3 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0_l~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0_l~3 .extended_lut = "off";
defparam \cal_pd0_l~3 .lut_mask = 64'h0101010101010101;
defparam \cal_pd0_l~3 .shared_arith = "off";

dffeas \cal_pd0_l[1] (
	.clk(clock),
	.d(\cal_pd0_l~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd0_l[0]~1_combout ),
	.q(\cal_pd0_l[1]~q ),
	.prn(vcc));
defparam \cal_pd0_l[1] .is_wysiwyg = "true";
defparam \cal_pd0_l[1] .power_up = "low";

cyclonev_lcell_comb \cal_pd0_l~2 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0_l~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0_l~2 .extended_lut = "off";
defparam \cal_pd0_l~2 .lut_mask = 64'h0101010101010101;
defparam \cal_pd0_l~2 .shared_arith = "off";

dffeas \cal_pd0_l[0] (
	.clk(clock),
	.d(\cal_pd0_l~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd0_l[0]~1_combout ),
	.q(\cal_pd0_l[0]~q ),
	.prn(vcc));
defparam \cal_pd0_l[0] .is_wysiwyg = "true";
defparam \cal_pd0_l[0] .power_up = "low";

cyclonev_lcell_comb \Add0~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd0[0]~q ),
	.datae(gnd),
	.dataf(!\cal_pd0_l[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~18_cout ),
	.shareout());
defparam \Add0~18 .extended_lut = "off";
defparam \Add0~18 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~18 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd0[1]~q ),
	.datae(gnd),
	.dataf(!\cal_pd0_l[1]~q ),
	.datag(gnd),
	.cin(\Add0~18_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd0[2]~q ),
	.datae(gnd),
	.dataf(!\cal_pd0_l[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd0~0 (
	.dataa(!\cal_pd0[0]~q ),
	.datab(!\cal_pd0[3]~q ),
	.datac(!\cal_pd0[2]~q ),
	.datad(!\cal_pd0[1]~q ),
	.datae(!\cal_inc[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0~0 .extended_lut = "off";
defparam \cal_pd0~0 .lut_mask = 64'h0001000000010000;
defparam \cal_pd0~0 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd0~3 (
	.dataa(!\cal_done[0]~q ),
	.datab(!\cal_pd0~0_combout ),
	.datac(!\cal_pd0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0~3 .extended_lut = "off";
defparam \cal_pd0~3 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \cal_pd0~3 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd0~6 (
	.dataa(!\cal_inc[0]~q ),
	.datab(!\cal_pd0~2_combout ),
	.datac(!\Add0~5_sumout ),
	.datad(!\cal_pd0~1_combout ),
	.datae(!\cal_pd0~3_combout ),
	.dataf(!\cal_pd0[1]~q ),
	.datag(!\cal_pd0[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0~6 .extended_lut = "on";
defparam \cal_pd0~6 .lut_mask = 64'h12123F0CEDED3F0C;
defparam \cal_pd0~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[1]~q ),
	.datad(!\cal_pd0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector24~0 .shared_arith = "off";

dffeas \cal_pd0[1] (
	.clk(clock),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd0[1]~q ),
	.prn(vcc));
defparam \cal_pd0[1] .is_wysiwyg = "true";
defparam \cal_pd0[1] .power_up = "low";

cyclonev_lcell_comb \Add6~1 (
	.dataa(!\cal_pd0[0]~q ),
	.datab(!\cal_pd0[2]~q ),
	.datac(!\cal_pd0[1]~q ),
	.datad(!\cal_inc[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add6~1 .extended_lut = "off";
defparam \Add6~1 .lut_mask = 64'h3693369336933693;
defparam \Add6~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd0[3]~q ),
	.datae(gnd),
	.dataf(!\cal_pd0_l[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd0~5 (
	.dataa(!\cal_pd0[2]~q ),
	.datab(!\Add6~1_combout ),
	.datac(!\Add0~13_sumout ),
	.datad(!\cal_pd0~1_combout ),
	.datae(!\cal_pd0~2_combout ),
	.dataf(!\cal_pd0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0~5 .extended_lut = "off";
defparam \cal_pd0~5 .lut_mask = 64'h555533330F0FFF00;
defparam \cal_pd0~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector23~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[2]~q ),
	.datad(!\cal_pd0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector23~0 .shared_arith = "off";

dffeas \cal_pd0[2] (
	.clk(clock),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd0[2]~q ),
	.prn(vcc));
defparam \cal_pd0[2] .is_wysiwyg = "true";
defparam \cal_pd0[2] .power_up = "low";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!\cal_pd0[0]~q ),
	.datab(!\cal_pd0[2]~q ),
	.datac(!\cal_pd0[1]~q ),
	.datad(!\cal_pd0_l[0]~q ),
	.datae(!\cal_pd0_l[1]~q ),
	.dataf(!\cal_pd0_l[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h8040080420100201;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector65~0 (
	.dataa(!\cal_pd0[3]~q ),
	.datab(!\cal_inc[0]~q ),
	.datac(!\cal_pd0_l[3]~q ),
	.datad(!\Equal4~0_combout ),
	.datae(!\cal_pd0~0_combout ),
	.dataf(!\cal_pd0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector65~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector65~0 .extended_lut = "off";
defparam \Selector65~0 .lut_mask = 64'h00000000FFDE0000;
defparam \Selector65~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector65~1 (
	.dataa(!\cal_done[0]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\WideOr8~0_combout ),
	.datad(!\Selector57~2_combout ),
	.datae(!\ignore_solid[0]~q ),
	.dataf(!\Selector65~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector65~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector65~1 .extended_lut = "off";
defparam \Selector65~1 .lut_mask = 64'hE000FFFFC000DDDD;
defparam \Selector65~1 .shared_arith = "off";

dffeas \ignore_solid[0] (
	.clk(clock),
	.d(\Selector65~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ignore_solid[0]~q ),
	.prn(vcc));
defparam \ignore_solid[0] .is_wysiwyg = "true";
defparam \ignore_solid[0] .power_up = "low";

dffeas \data_e0q[0] (
	.clk(clock),
	.d(\pd0_det|ff2~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e0q[0]~q ),
	.prn(vcc));
defparam \data_e0q[0] .is_wysiwyg = "true";
defparam \data_e0q[0] .power_up = "low";

dffeas \data_e1q[0] (
	.clk(clock),
	.d(\data_e0q[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e1q[0]~q ),
	.prn(vcc));
defparam \data_e1q[0] .is_wysiwyg = "true";
defparam \data_e1q[0] .power_up = "low";

cyclonev_lcell_comb \cal_pd0~1 (
	.dataa(!\pd_0_p[0]~q ),
	.datab(!\pd_0[0]~q ),
	.datac(!\pd_1_p[0]~q ),
	.datad(!\pd_1[0]~q ),
	.datae(!\ignore_solid[0]~q ),
	.dataf(!\data_e1q[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0~1 .extended_lut = "off";
defparam \cal_pd0~1 .lut_mask = 64'hF99FFFFF00000000;
defparam \cal_pd0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector61~0 (
	.dataa(!\cal_done[0]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\cal_inc[0]~q ),
	.datae(!\cal_pd0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector61~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector61~0 .extended_lut = "off";
defparam \Selector61~0 .lut_mask = 64'h22F200F022F200F0;
defparam \Selector61~0 .shared_arith = "off";

dffeas \cal_inc[0] (
	.clk(clock),
	.d(\Selector61~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_inc[0]~q ),
	.prn(vcc));
defparam \cal_inc[0] .is_wysiwyg = "true";
defparam \cal_inc[0] .power_up = "low";

cyclonev_lcell_comb \cal_pd0~2 (
	.dataa(!\cal_done[0]~q ),
	.datab(!\cal_pd0[3]~q ),
	.datac(!\cal_inc[0]~q ),
	.datad(!\cal_pd0_l[3]~q ),
	.datae(!\Equal4~0_combout ),
	.dataf(!\cal_pd0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0~2 .extended_lut = "off";
defparam \cal_pd0~2 .lut_mask = 64'hA0A0A0A0AAAAA2A8;
defparam \cal_pd0~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!\cal_done[0]~q ),
	.datab(!\cal_pd0[0]~q ),
	.datac(!\cal_pd0~0_combout ),
	.datad(!\cal_pd0~1_combout ),
	.datae(!\Add0~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h1131BB3B1131BB3B;
defparam \Selector25~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~1 (
	.dataa(!\cal_done[0]~q ),
	.datab(!\cal_pd0[0]~q ),
	.datac(!\cal_pd0~0_combout ),
	.datad(!\cal_pd0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~1 .extended_lut = "off";
defparam \Selector25~1 .lut_mask = 64'h113B113B113B113B;
defparam \Selector25~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~2 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[0]~q ),
	.datad(!\cal_pd0~2_combout ),
	.datae(!\Selector25~0_combout ),
	.dataf(!\Selector25~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~2 .extended_lut = "off";
defparam \Selector25~2 .lut_mask = 64'h083B3B3B08083B08;
defparam \Selector25~2 .shared_arith = "off";

dffeas \cal_pd0[0] (
	.clk(clock),
	.d(\Selector25~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd0[0]~q ),
	.prn(vcc));
defparam \cal_pd0[0] .is_wysiwyg = "true";
defparam \cal_pd0[0] .power_up = "low";

cyclonev_lcell_comb \Add6~0 (
	.dataa(!\cal_pd0[0]~q ),
	.datab(!\cal_pd0[3]~q ),
	.datac(!\cal_pd0[2]~q ),
	.datad(!\cal_pd0[1]~q ),
	.datae(!\cal_inc[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add6~0 .extended_lut = "off";
defparam \Add6~0 .lut_mask = 64'h3336933333369333;
defparam \Add6~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FFFF00000000;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd0~4 (
	.dataa(!\cal_pd0[3]~q ),
	.datab(!\Add6~0_combout ),
	.datac(!\Add0~1_sumout ),
	.datad(!\cal_pd0~1_combout ),
	.datae(!\cal_pd0~2_combout ),
	.dataf(!\cal_pd0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd0~4 .extended_lut = "off";
defparam \cal_pd0~4 .lut_mask = 64'h555533330F0FFF00;
defparam \cal_pd0~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector22~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd0[3]~q ),
	.datad(!\cal_pd0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector22~0 .extended_lut = "off";
defparam \Selector22~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector22~0 .shared_arith = "off";

dffeas \cal_pd0[3] (
	.clk(clock),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd0[3]~q ),
	.prn(vcc));
defparam \cal_pd0[3] .is_wysiwyg = "true";
defparam \cal_pd0[3] .power_up = "low";

cyclonev_lcell_comb \Selector57~0 (
	.dataa(!\cal_pd0[3]~q ),
	.datab(!\cal_inc[0]~q ),
	.datac(!\cal_pd0_l[3]~q ),
	.datad(!\Equal4~0_combout ),
	.datae(!\cal_pd0~0_combout ),
	.dataf(!\cal_pd0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector57~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector57~0 .extended_lut = "off";
defparam \Selector57~0 .lut_mask = 64'hCCCCCCCCFFDE0000;
defparam \Selector57~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector57~1 (
	.dataa(!\cal_done[0]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\Selector57~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector57~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector57~1 .extended_lut = "off";
defparam \Selector57~1 .lut_mask = 64'h7350735073507350;
defparam \Selector57~1 .shared_arith = "off";

dffeas \cal_done[0] (
	.clk(clock),
	.d(\Selector57~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_done[0]~q ),
	.prn(vcc));
defparam \cal_done[0] .is_wysiwyg = "true";
defparam \cal_done[0] .power_up = "low";

dffeas \ch_testbus0q[1] (
	.clk(clock),
	.d(out_narrow_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus0q[1]~q ),
	.prn(vcc));
defparam \ch_testbus0q[1] .is_wysiwyg = "true";
defparam \ch_testbus0q[1] .power_up = "low";

dffeas \ch_testbus1q[1] (
	.clk(clock),
	.d(\ch_testbus0q[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus1q[1]~q ),
	.prn(vcc));
defparam \ch_testbus1q[1] .is_wysiwyg = "true";
defparam \ch_testbus1q[1] .power_up = "low";

cyclonev_lcell_comb \pd_0~2 (
	.dataa(!\pd_0[1]~q ),
	.datab(!\ch_testbus1q[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_0~2 .extended_lut = "off";
defparam \pd_0~2 .lut_mask = 64'h4444444444444444;
defparam \pd_0~2 .shared_arith = "off";

dffeas \pd_0[1] (
	.clk(clock),
	.d(\pd_0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_0[1]~q ),
	.prn(vcc));
defparam \pd_0[1] .is_wysiwyg = "true";
defparam \pd_0[1] .power_up = "low";

dffeas \pd_0_p[1] (
	.clk(clock),
	.d(\pd_0[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_0_p[1]~q ),
	.prn(vcc));
defparam \pd_0_p[1] .is_wysiwyg = "true";
defparam \pd_0_p[1] .power_up = "low";

cyclonev_lcell_comb \pd_1~1 (
	.dataa(!\pd_1[1]~q ),
	.datab(!\ch_testbus1q[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_1~1 .extended_lut = "off";
defparam \pd_1~1 .lut_mask = 64'h1111111111111111;
defparam \pd_1~1 .shared_arith = "off";

dffeas \pd_1[1] (
	.clk(clock),
	.d(\pd_1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_1[1]~q ),
	.prn(vcc));
defparam \pd_1[1] .is_wysiwyg = "true";
defparam \pd_1[1] .power_up = "low";

dffeas \pd_1_p[1] (
	.clk(clock),
	.d(\pd_1[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_1_p[1]~q ),
	.prn(vcc));
defparam \pd_1_p[1] .is_wysiwyg = "true";
defparam \pd_1_p[1] .power_up = "low";

cyclonev_lcell_comb \cal_pd90_l~0 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90_l~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90_l~0 .extended_lut = "off";
defparam \cal_pd90_l~0 .lut_mask = 64'h0101010101010101;
defparam \cal_pd90_l~0 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd90_l[3]~1 (
	.dataa(!reset),
	.datab(!\cal_done[1]~q ),
	.datac(!\state.TEST_INPUT~q ),
	.datad(!\Selector56~3_combout ),
	.datae(!\cal_inc[1]~q ),
	.dataf(!\cal_pd90~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90_l[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90_l[3]~1 .extended_lut = "off";
defparam \cal_pd90_l[3]~1 .lut_mask = 64'hAAFEAAFAAAFAAAFA;
defparam \cal_pd90_l[3]~1 .shared_arith = "off";

dffeas \cal_pd90_l[3] (
	.clk(clock),
	.d(\cal_pd90_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd90_l[3]~1_combout ),
	.q(\cal_pd90_l[3]~q ),
	.prn(vcc));
defparam \cal_pd90_l[3] .is_wysiwyg = "true";
defparam \cal_pd90_l[3] .power_up = "low";

cyclonev_lcell_comb \cal_pd90~2 (
	.dataa(!\cal_done[1]~q ),
	.datab(!\cal_pd90[3]~q ),
	.datac(!\cal_inc[1]~q ),
	.datad(!\cal_pd90_l[3]~q ),
	.datae(!\Equal6~0_combout ),
	.dataf(!\cal_pd90~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90~2 .extended_lut = "off";
defparam \cal_pd90~2 .lut_mask = 64'hA0A0A0A0AAAAA2A8;
defparam \cal_pd90~2 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd90~0 (
	.dataa(!\cal_pd90[3]~q ),
	.datab(!\cal_pd90[2]~q ),
	.datac(!\cal_pd90[1]~q ),
	.datad(!\cal_pd90[0]~q ),
	.datae(!\cal_inc[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90~0 .extended_lut = "off";
defparam \cal_pd90~0 .lut_mask = 64'h0001000000010000;
defparam \cal_pd90~0 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd90_l~3 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90_l~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90_l~3 .extended_lut = "off";
defparam \cal_pd90_l~3 .lut_mask = 64'h0101010101010101;
defparam \cal_pd90_l~3 .shared_arith = "off";

dffeas \cal_pd90_l[1] (
	.clk(clock),
	.d(\cal_pd90_l~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd90_l[3]~1_combout ),
	.q(\cal_pd90_l[1]~q ),
	.prn(vcc));
defparam \cal_pd90_l[1] .is_wysiwyg = "true";
defparam \cal_pd90_l[1] .power_up = "low";

cyclonev_lcell_comb \cal_pd90_l~2 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90_l~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90_l~2 .extended_lut = "off";
defparam \cal_pd90_l~2 .lut_mask = 64'h0101010101010101;
defparam \cal_pd90_l~2 .shared_arith = "off";

dffeas \cal_pd90_l[0] (
	.clk(clock),
	.d(\cal_pd90_l~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd90_l[3]~1_combout ),
	.q(\cal_pd90_l[0]~q ),
	.prn(vcc));
defparam \cal_pd90_l[0] .is_wysiwyg = "true";
defparam \cal_pd90_l[0] .power_up = "low";

cyclonev_lcell_comb \Add1~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd90[0]~q ),
	.datae(gnd),
	.dataf(!\cal_pd90_l[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add1~18_cout ),
	.shareout());
defparam \Add1~18 .extended_lut = "off";
defparam \Add1~18 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~18 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd90[1]~q ),
	.datae(gnd),
	.dataf(!\cal_pd90_l[1]~q ),
	.datag(gnd),
	.cin(\Add1~18_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!\cal_done[1]~q ),
	.datab(!\cal_pd90[0]~q ),
	.datac(!\cal_pd90~0_combout ),
	.datad(!\cal_pd90~1_combout ),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'h1131BB3B1131BB3B;
defparam \Selector29~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~1 (
	.dataa(!\cal_done[1]~q ),
	.datab(!\cal_pd90[0]~q ),
	.datac(!\cal_pd90~0_combout ),
	.datad(!\cal_pd90~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~1 .extended_lut = "off";
defparam \Selector29~1 .lut_mask = 64'h113B113B113B113B;
defparam \Selector29~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~2 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[0]~q ),
	.datad(!\cal_pd90~2_combout ),
	.datae(!\Selector29~0_combout ),
	.dataf(!\Selector29~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~2 .extended_lut = "off";
defparam \Selector29~2 .lut_mask = 64'h083B3B3B08083B08;
defparam \Selector29~2 .shared_arith = "off";

dffeas \cal_pd90[0] (
	.clk(clock),
	.d(\Selector29~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd90[0]~q ),
	.prn(vcc));
defparam \cal_pd90[0] .is_wysiwyg = "true";
defparam \cal_pd90[0] .power_up = "low";

cyclonev_lcell_comb \cal_pd90_l~4 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90_l~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90_l~4 .extended_lut = "off";
defparam \cal_pd90_l~4 .lut_mask = 64'h0101010101010101;
defparam \cal_pd90_l~4 .shared_arith = "off";

dffeas \cal_pd90_l[2] (
	.clk(clock),
	.d(\cal_pd90_l~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd90_l[3]~1_combout ),
	.q(\cal_pd90_l[2]~q ),
	.prn(vcc));
defparam \cal_pd90_l[2] .is_wysiwyg = "true";
defparam \cal_pd90_l[2] .power_up = "low";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!\cal_pd90[2]~q ),
	.datab(!\cal_pd90[1]~q ),
	.datac(!\cal_pd90[0]~q ),
	.datad(!\cal_pd90_l[0]~q ),
	.datae(!\cal_pd90_l[1]~q ),
	.dataf(!\cal_pd90_l[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h8008200240041001;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector64~0 (
	.dataa(!\cal_pd90[3]~q ),
	.datab(!\cal_inc[1]~q ),
	.datac(!\cal_pd90_l[3]~q ),
	.datad(!\Equal6~0_combout ),
	.datae(!\cal_pd90~0_combout ),
	.dataf(!\cal_pd90~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector64~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector64~0 .extended_lut = "off";
defparam \Selector64~0 .lut_mask = 64'h00000000FFDE0000;
defparam \Selector64~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector64~1 (
	.dataa(!\cal_done[1]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\WideOr8~0_combout ),
	.datad(!\Selector57~2_combout ),
	.datae(!\ignore_solid[1]~q ),
	.dataf(!\Selector64~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector64~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector64~1 .extended_lut = "off";
defparam \Selector64~1 .lut_mask = 64'hE000FFFFC000DDDD;
defparam \Selector64~1 .shared_arith = "off";

dffeas \ignore_solid[1] (
	.clk(clock),
	.d(\Selector64~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ignore_solid[1]~q ),
	.prn(vcc));
defparam \ignore_solid[1] .is_wysiwyg = "true";
defparam \ignore_solid[1] .power_up = "low";

dffeas \data_e0q[1] (
	.clk(clock),
	.d(\pd90_det|ff2~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e0q[1]~q ),
	.prn(vcc));
defparam \data_e0q[1] .is_wysiwyg = "true";
defparam \data_e0q[1] .power_up = "low";

dffeas \data_e1q[1] (
	.clk(clock),
	.d(\data_e0q[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e1q[1]~q ),
	.prn(vcc));
defparam \data_e1q[1] .is_wysiwyg = "true";
defparam \data_e1q[1] .power_up = "low";

cyclonev_lcell_comb \cal_pd90~1 (
	.dataa(!\pd_0_p[1]~q ),
	.datab(!\pd_0[1]~q ),
	.datac(!\pd_1_p[1]~q ),
	.datad(!\pd_1[1]~q ),
	.datae(!\ignore_solid[1]~q ),
	.dataf(!\data_e1q[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90~1 .extended_lut = "off";
defparam \cal_pd90~1 .lut_mask = 64'hF99FFFFF00000000;
defparam \cal_pd90~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector60~0 (
	.dataa(!\cal_done[1]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\cal_inc[1]~q ),
	.datae(!\cal_pd90~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector60~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector60~0 .extended_lut = "off";
defparam \Selector60~0 .lut_mask = 64'h22F200F022F200F0;
defparam \Selector60~0 .shared_arith = "off";

dffeas \cal_inc[1] (
	.clk(clock),
	.d(\Selector60~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_inc[1]~q ),
	.prn(vcc));
defparam \cal_inc[1] .is_wysiwyg = "true";
defparam \cal_inc[1] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd90[2]~q ),
	.datae(gnd),
	.dataf(!\cal_pd90_l[2]~q ),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd90~3 (
	.dataa(!\cal_done[1]~q ),
	.datab(!\cal_pd90~0_combout ),
	.datac(!\cal_pd90~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90~3 .extended_lut = "off";
defparam \cal_pd90~3 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \cal_pd90~3 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd90~6 (
	.dataa(!\cal_inc[1]~q ),
	.datab(!\cal_pd90~2_combout ),
	.datac(!\Add1~13_sumout ),
	.datad(!\cal_pd90~1_combout ),
	.datae(!\cal_pd90~3_combout ),
	.dataf(!\cal_pd90[1]~q ),
	.datag(!\cal_pd90[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90~6 .extended_lut = "on";
defparam \cal_pd90~6 .lut_mask = 64'h12123F0CEDED3F0C;
defparam \cal_pd90~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[1]~q ),
	.datad(!\cal_pd90~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector28~0 .shared_arith = "off";

dffeas \cal_pd90[1] (
	.clk(clock),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd90[1]~q ),
	.prn(vcc));
defparam \cal_pd90[1] .is_wysiwyg = "true";
defparam \cal_pd90[1] .power_up = "low";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!\cal_pd90[2]~q ),
	.datab(!\cal_pd90[1]~q ),
	.datac(!\cal_pd90[0]~q ),
	.datad(!\cal_inc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h5695569556955695;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd90[3]~q ),
	.datae(gnd),
	.dataf(!\cal_pd90_l[3]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd90~5 (
	.dataa(!\cal_pd90[2]~q ),
	.datab(!\Add7~1_combout ),
	.datac(!\Add1~9_sumout ),
	.datad(!\cal_pd90~1_combout ),
	.datae(!\cal_pd90~2_combout ),
	.dataf(!\cal_pd90~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90~5 .extended_lut = "off";
defparam \cal_pd90~5 .lut_mask = 64'h555533330F0FFF00;
defparam \cal_pd90~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[2]~q ),
	.datad(!\cal_pd90~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector27~0 .shared_arith = "off";

dffeas \cal_pd90[2] (
	.clk(clock),
	.d(\Selector27~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd90[2]~q ),
	.prn(vcc));
defparam \cal_pd90[2] .is_wysiwyg = "true";
defparam \cal_pd90[2] .power_up = "low";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!\cal_pd90[3]~q ),
	.datab(!\cal_pd90[2]~q ),
	.datac(!\cal_pd90[1]~q ),
	.datad(!\cal_pd90[0]~q ),
	.datae(!\cal_inc[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h5556955555569555;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FFFF00000000;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd90~4 (
	.dataa(!\cal_pd90[3]~q ),
	.datab(!\Add7~0_combout ),
	.datac(!\Add1~1_sumout ),
	.datad(!\cal_pd90~1_combout ),
	.datae(!\cal_pd90~2_combout ),
	.dataf(!\cal_pd90~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd90~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd90~4 .extended_lut = "off";
defparam \cal_pd90~4 .lut_mask = 64'h555533330F0FFF00;
defparam \cal_pd90~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd90[3]~q ),
	.datad(!\cal_pd90~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector26~0 .shared_arith = "off";

dffeas \cal_pd90[3] (
	.clk(clock),
	.d(\Selector26~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd90[3]~q ),
	.prn(vcc));
defparam \cal_pd90[3] .is_wysiwyg = "true";
defparam \cal_pd90[3] .power_up = "low";

cyclonev_lcell_comb \Selector56~1 (
	.dataa(!\cal_pd90[3]~q ),
	.datab(!\cal_inc[1]~q ),
	.datac(!\cal_pd90_l[3]~q ),
	.datad(!\Equal6~0_combout ),
	.datae(!\cal_pd90~0_combout ),
	.dataf(!\cal_pd90~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector56~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector56~1 .extended_lut = "off";
defparam \Selector56~1 .lut_mask = 64'hCCCCCCCCFFDE0000;
defparam \Selector56~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector56~2 (
	.dataa(!\cal_done[1]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\Selector56~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector56~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector56~2 .extended_lut = "off";
defparam \Selector56~2 .lut_mask = 64'h7350735073507350;
defparam \Selector56~2 .shared_arith = "off";

dffeas \cal_done[1] (
	.clk(clock),
	.d(\Selector56~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_done[1]~q ),
	.prn(vcc));
defparam \cal_done[1] .is_wysiwyg = "true";
defparam \cal_done[1] .power_up = "low";

dffeas \ch_testbus0q[2] (
	.clk(clock),
	.d(out_narrow_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus0q[2]~q ),
	.prn(vcc));
defparam \ch_testbus0q[2] .is_wysiwyg = "true";
defparam \ch_testbus0q[2] .power_up = "low";

dffeas \ch_testbus1q[2] (
	.clk(clock),
	.d(\ch_testbus0q[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus1q[2]~q ),
	.prn(vcc));
defparam \ch_testbus1q[2] .is_wysiwyg = "true";
defparam \ch_testbus1q[2] .power_up = "low";

cyclonev_lcell_comb \pd_0~3 (
	.dataa(!\pd_0[2]~q ),
	.datab(!\ch_testbus1q[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_0~3 .extended_lut = "off";
defparam \pd_0~3 .lut_mask = 64'h4444444444444444;
defparam \pd_0~3 .shared_arith = "off";

dffeas \pd_0[2] (
	.clk(clock),
	.d(\pd_0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_0[2]~q ),
	.prn(vcc));
defparam \pd_0[2] .is_wysiwyg = "true";
defparam \pd_0[2] .power_up = "low";

dffeas \pd_0_p[2] (
	.clk(clock),
	.d(\pd_0[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_0_p[2]~q ),
	.prn(vcc));
defparam \pd_0_p[2] .is_wysiwyg = "true";
defparam \pd_0_p[2] .power_up = "low";

cyclonev_lcell_comb \pd_1~2 (
	.dataa(!\pd_1[2]~q ),
	.datab(!\ch_testbus1q[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_1~2 .extended_lut = "off";
defparam \pd_1~2 .lut_mask = 64'h1111111111111111;
defparam \pd_1~2 .shared_arith = "off";

dffeas \pd_1[2] (
	.clk(clock),
	.d(\pd_1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_1[2]~q ),
	.prn(vcc));
defparam \pd_1[2] .is_wysiwyg = "true";
defparam \pd_1[2] .power_up = "low";

dffeas \pd_1_p[2] (
	.clk(clock),
	.d(\pd_1[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_1_p[2]~q ),
	.prn(vcc));
defparam \pd_1_p[2] .is_wysiwyg = "true";
defparam \pd_1_p[2] .power_up = "low";

cyclonev_lcell_comb \cal_pd180_l~0 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180_l~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180_l~0 .extended_lut = "off";
defparam \cal_pd180_l~0 .lut_mask = 64'h0101010101010101;
defparam \cal_pd180_l~0 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd180_l[3]~1 (
	.dataa(!reset),
	.datab(!\cal_done[2]~q ),
	.datac(!\state.TEST_INPUT~q ),
	.datad(!\Selector56~3_combout ),
	.datae(!\cal_inc[2]~q ),
	.dataf(!\cal_pd180~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180_l[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180_l[3]~1 .extended_lut = "off";
defparam \cal_pd180_l[3]~1 .lut_mask = 64'hAAFEAAFAAAFAAAFA;
defparam \cal_pd180_l[3]~1 .shared_arith = "off";

dffeas \cal_pd180_l[3] (
	.clk(clock),
	.d(\cal_pd180_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd180_l[3]~1_combout ),
	.q(\cal_pd180_l[3]~q ),
	.prn(vcc));
defparam \cal_pd180_l[3] .is_wysiwyg = "true";
defparam \cal_pd180_l[3] .power_up = "low";

cyclonev_lcell_comb \cal_pd180~2 (
	.dataa(!\cal_done[2]~q ),
	.datab(!\cal_pd180[3]~q ),
	.datac(!\cal_inc[2]~q ),
	.datad(!\cal_pd180_l[3]~q ),
	.datae(!\Equal8~0_combout ),
	.dataf(!\cal_pd180~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180~2 .extended_lut = "off";
defparam \cal_pd180~2 .lut_mask = 64'hA0A0A0A0AAAAA2A8;
defparam \cal_pd180~2 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd180~0 (
	.dataa(!\cal_pd180[3]~q ),
	.datab(!\cal_pd180[2]~q ),
	.datac(!\cal_pd180[1]~q ),
	.datad(!\cal_pd180[0]~q ),
	.datae(!\cal_inc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180~0 .extended_lut = "off";
defparam \cal_pd180~0 .lut_mask = 64'h0001000000010000;
defparam \cal_pd180~0 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd180_l~3 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180_l~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180_l~3 .extended_lut = "off";
defparam \cal_pd180_l~3 .lut_mask = 64'h0101010101010101;
defparam \cal_pd180_l~3 .shared_arith = "off";

dffeas \cal_pd180_l[1] (
	.clk(clock),
	.d(\cal_pd180_l~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd180_l[3]~1_combout ),
	.q(\cal_pd180_l[1]~q ),
	.prn(vcc));
defparam \cal_pd180_l[1] .is_wysiwyg = "true";
defparam \cal_pd180_l[1] .power_up = "low";

cyclonev_lcell_comb \cal_pd180_l~2 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180_l~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180_l~2 .extended_lut = "off";
defparam \cal_pd180_l~2 .lut_mask = 64'h0101010101010101;
defparam \cal_pd180_l~2 .shared_arith = "off";

dffeas \cal_pd180_l[0] (
	.clk(clock),
	.d(\cal_pd180_l~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd180_l[3]~1_combout ),
	.q(\cal_pd180_l[0]~q ),
	.prn(vcc));
defparam \cal_pd180_l[0] .is_wysiwyg = "true";
defparam \cal_pd180_l[0] .power_up = "low";

cyclonev_lcell_comb \Add2~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd180[0]~q ),
	.datae(gnd),
	.dataf(!\cal_pd180_l[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add2~18_cout ),
	.shareout());
defparam \Add2~18 .extended_lut = "off";
defparam \Add2~18 .lut_mask = 64'h0000FF00000000FF;
defparam \Add2~18 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd180[1]~q ),
	.datae(gnd),
	.dataf(!\cal_pd180_l[1]~q ),
	.datag(gnd),
	.cin(\Add2~18_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector33~0 (
	.dataa(!\cal_done[2]~q ),
	.datab(!\cal_pd180[0]~q ),
	.datac(!\cal_pd180~0_combout ),
	.datad(!\cal_pd180~1_combout ),
	.datae(!\Add2~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~0 .extended_lut = "off";
defparam \Selector33~0 .lut_mask = 64'h1131BB3B1131BB3B;
defparam \Selector33~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector33~1 (
	.dataa(!\cal_done[2]~q ),
	.datab(!\cal_pd180[0]~q ),
	.datac(!\cal_pd180~0_combout ),
	.datad(!\cal_pd180~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~1 .extended_lut = "off";
defparam \Selector33~1 .lut_mask = 64'h113B113B113B113B;
defparam \Selector33~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector33~2 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[0]~q ),
	.datad(!\cal_pd180~2_combout ),
	.datae(!\Selector33~0_combout ),
	.dataf(!\Selector33~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~2 .extended_lut = "off";
defparam \Selector33~2 .lut_mask = 64'h083B3B3B08083B08;
defparam \Selector33~2 .shared_arith = "off";

dffeas \cal_pd180[0] (
	.clk(clock),
	.d(\Selector33~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd180[0]~q ),
	.prn(vcc));
defparam \cal_pd180[0] .is_wysiwyg = "true";
defparam \cal_pd180[0] .power_up = "low";

cyclonev_lcell_comb \cal_pd180_l~4 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180_l~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180_l~4 .extended_lut = "off";
defparam \cal_pd180_l~4 .lut_mask = 64'h0101010101010101;
defparam \cal_pd180_l~4 .shared_arith = "off";

dffeas \cal_pd180_l[2] (
	.clk(clock),
	.d(\cal_pd180_l~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd180_l[3]~1_combout ),
	.q(\cal_pd180_l[2]~q ),
	.prn(vcc));
defparam \cal_pd180_l[2] .is_wysiwyg = "true";
defparam \cal_pd180_l[2] .power_up = "low";

cyclonev_lcell_comb \Equal8~0 (
	.dataa(!\cal_pd180[2]~q ),
	.datab(!\cal_pd180[1]~q ),
	.datac(!\cal_pd180[0]~q ),
	.datad(!\cal_pd180_l[0]~q ),
	.datae(!\cal_pd180_l[1]~q ),
	.dataf(!\cal_pd180_l[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal8~0 .extended_lut = "off";
defparam \Equal8~0 .lut_mask = 64'h8008200240041001;
defparam \Equal8~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector63~0 (
	.dataa(!\cal_pd180[3]~q ),
	.datab(!\cal_inc[2]~q ),
	.datac(!\cal_pd180_l[3]~q ),
	.datad(!\Equal8~0_combout ),
	.datae(!\cal_pd180~0_combout ),
	.dataf(!\cal_pd180~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector63~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector63~0 .extended_lut = "off";
defparam \Selector63~0 .lut_mask = 64'h00000000FFDE0000;
defparam \Selector63~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector63~1 (
	.dataa(!\cal_done[2]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\WideOr8~0_combout ),
	.datad(!\Selector57~2_combout ),
	.datae(!\ignore_solid[2]~q ),
	.dataf(!\Selector63~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector63~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector63~1 .extended_lut = "off";
defparam \Selector63~1 .lut_mask = 64'hE000FFFFC000DDDD;
defparam \Selector63~1 .shared_arith = "off";

dffeas \ignore_solid[2] (
	.clk(clock),
	.d(\Selector63~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ignore_solid[2]~q ),
	.prn(vcc));
defparam \ignore_solid[2] .is_wysiwyg = "true";
defparam \ignore_solid[2] .power_up = "low";

dffeas \data_e0q[2] (
	.clk(clock),
	.d(\pd180_det|ff2~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e0q[2]~q ),
	.prn(vcc));
defparam \data_e0q[2] .is_wysiwyg = "true";
defparam \data_e0q[2] .power_up = "low";

dffeas \data_e1q[2] (
	.clk(clock),
	.d(\data_e0q[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e1q[2]~q ),
	.prn(vcc));
defparam \data_e1q[2] .is_wysiwyg = "true";
defparam \data_e1q[2] .power_up = "low";

cyclonev_lcell_comb \cal_pd180~1 (
	.dataa(!\pd_0_p[2]~q ),
	.datab(!\pd_0[2]~q ),
	.datac(!\pd_1_p[2]~q ),
	.datad(!\pd_1[2]~q ),
	.datae(!\ignore_solid[2]~q ),
	.dataf(!\data_e1q[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180~1 .extended_lut = "off";
defparam \cal_pd180~1 .lut_mask = 64'hF99FFFFF00000000;
defparam \cal_pd180~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector59~0 (
	.dataa(!\cal_done[2]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\cal_inc[2]~q ),
	.datae(!\cal_pd180~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector59~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector59~0 .extended_lut = "off";
defparam \Selector59~0 .lut_mask = 64'h22F200F022F200F0;
defparam \Selector59~0 .shared_arith = "off";

dffeas \cal_inc[2] (
	.clk(clock),
	.d(\Selector59~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_inc[2]~q ),
	.prn(vcc));
defparam \cal_inc[2] .is_wysiwyg = "true";
defparam \cal_inc[2] .power_up = "low";

cyclonev_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd180[2]~q ),
	.datae(gnd),
	.dataf(!\cal_pd180_l[2]~q ),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd180~3 (
	.dataa(!\cal_done[2]~q ),
	.datab(!\cal_pd180~0_combout ),
	.datac(!\cal_pd180~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180~3 .extended_lut = "off";
defparam \cal_pd180~3 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \cal_pd180~3 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd180~6 (
	.dataa(!\cal_inc[2]~q ),
	.datab(!\cal_pd180~2_combout ),
	.datac(!\Add2~13_sumout ),
	.datad(!\cal_pd180~1_combout ),
	.datae(!\cal_pd180~3_combout ),
	.dataf(!\cal_pd180[1]~q ),
	.datag(!\cal_pd180[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180~6 .extended_lut = "on";
defparam \cal_pd180~6 .lut_mask = 64'h12123F0CEDED3F0C;
defparam \cal_pd180~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector32~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[1]~q ),
	.datad(!\cal_pd180~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~0 .extended_lut = "off";
defparam \Selector32~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector32~0 .shared_arith = "off";

dffeas \cal_pd180[1] (
	.clk(clock),
	.d(\Selector32~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd180[1]~q ),
	.prn(vcc));
defparam \cal_pd180[1] .is_wysiwyg = "true";
defparam \cal_pd180[1] .power_up = "low";

cyclonev_lcell_comb \Add8~1 (
	.dataa(!\cal_pd180[2]~q ),
	.datab(!\cal_pd180[1]~q ),
	.datac(!\cal_pd180[0]~q ),
	.datad(!\cal_inc[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add8~1 .extended_lut = "off";
defparam \Add8~1 .lut_mask = 64'h5695569556955695;
defparam \Add8~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd180[3]~q ),
	.datae(gnd),
	.dataf(!\cal_pd180_l[3]~q ),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd180~5 (
	.dataa(!\cal_pd180[2]~q ),
	.datab(!\Add8~1_combout ),
	.datac(!\Add2~9_sumout ),
	.datad(!\cal_pd180~1_combout ),
	.datae(!\cal_pd180~2_combout ),
	.dataf(!\cal_pd180~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180~5 .extended_lut = "off";
defparam \cal_pd180~5 .lut_mask = 64'h555533330F0FFF00;
defparam \cal_pd180~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector31~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[2]~q ),
	.datad(!\cal_pd180~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector31~0 .extended_lut = "off";
defparam \Selector31~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector31~0 .shared_arith = "off";

dffeas \cal_pd180[2] (
	.clk(clock),
	.d(\Selector31~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd180[2]~q ),
	.prn(vcc));
defparam \cal_pd180[2] .is_wysiwyg = "true";
defparam \cal_pd180[2] .power_up = "low";

cyclonev_lcell_comb \Add8~0 (
	.dataa(!\cal_pd180[3]~q ),
	.datab(!\cal_pd180[2]~q ),
	.datac(!\cal_pd180[1]~q ),
	.datad(!\cal_pd180[0]~q ),
	.datae(!\cal_inc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add8~0 .extended_lut = "off";
defparam \Add8~0 .lut_mask = 64'h5556955555569555;
defparam \Add8~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FFFF00000000;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd180~4 (
	.dataa(!\cal_pd180[3]~q ),
	.datab(!\Add8~0_combout ),
	.datac(!\Add2~1_sumout ),
	.datad(!\cal_pd180~1_combout ),
	.datae(!\cal_pd180~2_combout ),
	.dataf(!\cal_pd180~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd180~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd180~4 .extended_lut = "off";
defparam \cal_pd180~4 .lut_mask = 64'h555533330F0FFF00;
defparam \cal_pd180~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector30~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd180[3]~q ),
	.datad(!\cal_pd180~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector30~0 .extended_lut = "off";
defparam \Selector30~0 .lut_mask = 64'h083B083B083B083B;
defparam \Selector30~0 .shared_arith = "off";

dffeas \cal_pd180[3] (
	.clk(clock),
	.d(\Selector30~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd180[3]~q ),
	.prn(vcc));
defparam \cal_pd180[3] .is_wysiwyg = "true";
defparam \cal_pd180[3] .power_up = "low";

cyclonev_lcell_comb \Selector55~0 (
	.dataa(!\cal_pd180[3]~q ),
	.datab(!\cal_inc[2]~q ),
	.datac(!\cal_pd180_l[3]~q ),
	.datad(!\Equal8~0_combout ),
	.datae(!\cal_pd180~0_combout ),
	.dataf(!\cal_pd180~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector55~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector55~0 .extended_lut = "off";
defparam \Selector55~0 .lut_mask = 64'hCCCCCCCCFFDE0000;
defparam \Selector55~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector55~1 (
	.dataa(!\cal_done[2]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\Selector55~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector55~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector55~1 .extended_lut = "off";
defparam \Selector55~1 .lut_mask = 64'h7350735073507350;
defparam \Selector55~1 .shared_arith = "off";

dffeas \cal_done[2] (
	.clk(clock),
	.d(\Selector55~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_done[2]~q ),
	.prn(vcc));
defparam \cal_done[2] .is_wysiwyg = "true";
defparam \cal_done[2] .power_up = "low";

dffeas \ch_testbus0q[3] (
	.clk(clock),
	.d(out_narrow_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus0q[3]~q ),
	.prn(vcc));
defparam \ch_testbus0q[3] .is_wysiwyg = "true";
defparam \ch_testbus0q[3] .power_up = "low";

dffeas \ch_testbus1q[3] (
	.clk(clock),
	.d(\ch_testbus0q[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ch_testbus1q[3]~q ),
	.prn(vcc));
defparam \ch_testbus1q[3] .is_wysiwyg = "true";
defparam \ch_testbus1q[3] .power_up = "low";

cyclonev_lcell_comb \pd_0~4 (
	.dataa(!\pd_0[3]~q ),
	.datab(!\ch_testbus1q[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_0~4 .extended_lut = "off";
defparam \pd_0~4 .lut_mask = 64'h4444444444444444;
defparam \pd_0~4 .shared_arith = "off";

dffeas \pd_0[3] (
	.clk(clock),
	.d(\pd_0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_0[3]~q ),
	.prn(vcc));
defparam \pd_0[3] .is_wysiwyg = "true";
defparam \pd_0[3] .power_up = "low";

dffeas \pd_0_p[3] (
	.clk(clock),
	.d(\pd_0[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_0_p[3]~q ),
	.prn(vcc));
defparam \pd_0_p[3] .is_wysiwyg = "true";
defparam \pd_0_p[3] .power_up = "low";

cyclonev_lcell_comb \pd_1~3 (
	.dataa(!\pd_1[3]~q ),
	.datab(!\ch_testbus1q[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_1~3 .extended_lut = "off";
defparam \pd_1~3 .lut_mask = 64'h1111111111111111;
defparam \pd_1~3 .shared_arith = "off";

dffeas \pd_1[3] (
	.clk(clock),
	.d(\pd_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\state.SAMPLE_TB~q ),
	.ena(\pd_0[0]~1_combout ),
	.q(\pd_1[3]~q ),
	.prn(vcc));
defparam \pd_1[3] .is_wysiwyg = "true";
defparam \pd_1[3] .power_up = "low";

dffeas \pd_1_p[3] (
	.clk(clock),
	.d(\pd_1[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pd_0_p[0]~1_combout ),
	.q(\pd_1_p[3]~q ),
	.prn(vcc));
defparam \pd_1_p[3] .is_wysiwyg = "true";
defparam \pd_1_p[3] .power_up = "low";

cyclonev_lcell_comb \Selector58~0 (
	.dataa(!\cal_done[3]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\cal_inc[3]~q ),
	.datae(!\edges[3]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector58~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector58~0 .extended_lut = "off";
defparam \Selector58~0 .lut_mask = 64'h22F200F022F200F0;
defparam \Selector58~0 .shared_arith = "off";

dffeas \cal_inc[3] (
	.clk(clock),
	.d(\Selector58~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_inc[3]~q ),
	.prn(vcc));
defparam \cal_inc[3] .is_wysiwyg = "true";
defparam \cal_inc[3] .power_up = "low";

cyclonev_lcell_comb \cal_pd270_l~0 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd270[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270_l~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270_l~0 .extended_lut = "off";
defparam \cal_pd270_l~0 .lut_mask = 64'h0101010101010101;
defparam \cal_pd270_l~0 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd270_l[1]~1 (
	.dataa(!reset),
	.datab(!\cal_done[3]~q ),
	.datac(!\state.TEST_INPUT~q ),
	.datad(!\Selector56~3_combout ),
	.datae(!\cal_inc[3]~q ),
	.dataf(!\edges[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270_l[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270_l[1]~1 .extended_lut = "off";
defparam \cal_pd270_l[1]~1 .lut_mask = 64'hAAFEAAFAAAFAAAFA;
defparam \cal_pd270_l[1]~1 .shared_arith = "off";

dffeas \cal_pd270_l[3] (
	.clk(clock),
	.d(\cal_pd270_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd270_l[1]~1_combout ),
	.q(\cal_pd270_l[3]~q ),
	.prn(vcc));
defparam \cal_pd270_l[3] .is_wysiwyg = "true";
defparam \cal_pd270_l[3] .power_up = "low";

cyclonev_lcell_comb \Add9~1 (
	.dataa(!\cal_pd270[0]~q ),
	.datab(!\cal_pd270[2]~q ),
	.datac(!\cal_pd270[1]~q ),
	.datad(!\cal_inc[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add9~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add9~1 .extended_lut = "off";
defparam \Add9~1 .lut_mask = 64'h3693369336933693;
defparam \Add9~1 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd270_l~4 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd270[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270_l~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270_l~4 .extended_lut = "off";
defparam \cal_pd270_l~4 .lut_mask = 64'h0101010101010101;
defparam \cal_pd270_l~4 .shared_arith = "off";

dffeas \cal_pd270_l[2] (
	.clk(clock),
	.d(\cal_pd270_l~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd270_l[1]~1_combout ),
	.q(\cal_pd270_l[2]~q ),
	.prn(vcc));
defparam \cal_pd270_l[2] .is_wysiwyg = "true";
defparam \cal_pd270_l[2] .power_up = "low";

cyclonev_lcell_comb \cal_pd270_l~3 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd270[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270_l~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270_l~3 .extended_lut = "off";
defparam \cal_pd270_l~3 .lut_mask = 64'h0101010101010101;
defparam \cal_pd270_l~3 .shared_arith = "off";

dffeas \cal_pd270_l[1] (
	.clk(clock),
	.d(\cal_pd270_l~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd270_l[1]~1_combout ),
	.q(\cal_pd270_l[1]~q ),
	.prn(vcc));
defparam \cal_pd270_l[1] .is_wysiwyg = "true";
defparam \cal_pd270_l[1] .power_up = "low";

cyclonev_lcell_comb \cal_pd270_l~2 (
	.dataa(!reset),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd270[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270_l~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270_l~2 .extended_lut = "off";
defparam \cal_pd270_l~2 .lut_mask = 64'h0101010101010101;
defparam \cal_pd270_l~2 .shared_arith = "off";

dffeas \cal_pd270_l[0] (
	.clk(clock),
	.d(\cal_pd270_l~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cal_pd270_l[1]~1_combout ),
	.q(\cal_pd270_l[0]~q ),
	.prn(vcc));
defparam \cal_pd270_l[0] .is_wysiwyg = "true";
defparam \cal_pd270_l[0] .power_up = "low";

cyclonev_lcell_comb \Add3~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd270[0]~q ),
	.datae(gnd),
	.dataf(!\cal_pd270_l[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add3~18_cout ),
	.shareout());
defparam \Add3~18 .extended_lut = "off";
defparam \Add3~18 .lut_mask = 64'h0000FF00000000FF;
defparam \Add3~18 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd270[1]~q ),
	.datae(gnd),
	.dataf(!\cal_pd270_l[1]~q ),
	.datag(gnd),
	.cin(\Add3~18_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd270[2]~q ),
	.datae(gnd),
	.dataf(!\cal_pd270_l[2]~q ),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add3~13 .shared_arith = "off";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cal_pd270[3]~q ),
	.datae(gnd),
	.dataf(!\cal_pd270_l[3]~q ),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add3~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector35~0 (
	.dataa(!\cal_done[3]~q ),
	.datab(!\cal_pd270[2]~q ),
	.datac(!\cal_pd270~0_combout ),
	.datad(!\cal_pd270~2_combout ),
	.datae(!\Add9~1_combout ),
	.dataf(!\Add3~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~0 .extended_lut = "off";
defparam \Selector35~0 .lut_mask = 64'hCEF0C4F0CE00C400;
defparam \Selector35~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector35~1 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd270[2]~q ),
	.datad(!\Selector35~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~1 .extended_lut = "off";
defparam \Selector35~1 .lut_mask = 64'h3B083B083B083B08;
defparam \Selector35~1 .shared_arith = "off";

dffeas \cal_pd270[2] (
	.clk(clock),
	.d(\Selector35~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd270[2]~q ),
	.prn(vcc));
defparam \cal_pd270[2] .is_wysiwyg = "true";
defparam \cal_pd270[2] .power_up = "low";

cyclonev_lcell_comb \cal_pd270~1 (
	.dataa(!\cal_pd270[0]~q ),
	.datab(!\cal_pd270[3]~q ),
	.datac(!\cal_pd270[2]~q ),
	.datad(!\cal_pd270[1]~q ),
	.datae(!\cal_inc[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270~1 .extended_lut = "off";
defparam \cal_pd270~1 .lut_mask = 64'h0001000000010000;
defparam \cal_pd270~1 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd270~2 (
	.dataa(!\cal_done[3]~q ),
	.datab(!\edges[3]~0_combout ),
	.datac(!\cal_pd270~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270~2 .extended_lut = "off";
defparam \cal_pd270~2 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \cal_pd270~2 .shared_arith = "off";

cyclonev_lcell_comb \Add9~2 (
	.dataa(!\cal_pd270[0]~q ),
	.datab(!\cal_pd270[1]~q ),
	.datac(!\cal_inc[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add9~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add9~2 .extended_lut = "off";
defparam \Add9~2 .lut_mask = 64'h6969696969696969;
defparam \Add9~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector36~0 (
	.dataa(!\cal_done[3]~q ),
	.datab(!\cal_pd270[1]~q ),
	.datac(!\cal_pd270~0_combout ),
	.datad(!\cal_pd270~2_combout ),
	.datae(!\Add9~2_combout ),
	.dataf(!\Add3~13_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~0 .extended_lut = "off";
defparam \Selector36~0 .lut_mask = 64'hCEF0C4F0CE00C400;
defparam \Selector36~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector36~1 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd270[1]~q ),
	.datad(!\Selector36~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~1 .extended_lut = "off";
defparam \Selector36~1 .lut_mask = 64'h3B083B083B083B08;
defparam \Selector36~1 .shared_arith = "off";

dffeas \cal_pd270[1] (
	.clk(clock),
	.d(\Selector36~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd270[1]~q ),
	.prn(vcc));
defparam \cal_pd270[1] .is_wysiwyg = "true";
defparam \cal_pd270[1] .power_up = "low";

cyclonev_lcell_comb \Selector37~0 (
	.dataa(!\cal_pd270~0_combout ),
	.datab(!\cal_pd270[0]~q ),
	.datac(!\Add3~1_sumout ),
	.datad(!\state.TEST_INPUT~q ),
	.datae(!\cal_pd270~2_combout ),
	.dataf(!\state.CH_WAIT~q ),
	.datag(!\cal_done[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector37~0 .extended_lut = "on";
defparam \Selector37~0 .lut_mask = 64'h3363335F0063005F;
defparam \Selector37~0 .shared_arith = "off";

dffeas \cal_pd270[0] (
	.clk(clock),
	.d(\Selector37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd270[0]~q ),
	.prn(vcc));
defparam \cal_pd270[0] .is_wysiwyg = "true";
defparam \cal_pd270[0] .power_up = "low";

cyclonev_lcell_comb \Equal10~0 (
	.dataa(!\cal_pd270[0]~q ),
	.datab(!\cal_pd270[2]~q ),
	.datac(!\cal_pd270[1]~q ),
	.datad(!\cal_pd270_l[0]~q ),
	.datae(!\cal_pd270_l[1]~q ),
	.dataf(!\cal_pd270_l[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal10~0 .extended_lut = "off";
defparam \Equal10~0 .lut_mask = 64'h8040080420100201;
defparam \Equal10~0 .shared_arith = "off";

cyclonev_lcell_comb \cal_pd270~0 (
	.dataa(!\cal_pd270[3]~q ),
	.datab(!\cal_inc[3]~q ),
	.datac(!\cal_pd270_l[3]~q ),
	.datad(!\edges[3]~0_combout ),
	.datae(!\Equal10~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_pd270~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cal_pd270~0 .extended_lut = "off";
defparam \cal_pd270~0 .lut_mask = 64'hCCFFCCDECCFFCCDE;
defparam \cal_pd270~0 .shared_arith = "off";

cyclonev_lcell_comb \Add9~0 (
	.dataa(!\cal_pd270[0]~q ),
	.datab(!\cal_pd270[3]~q ),
	.datac(!\cal_pd270[2]~q ),
	.datad(!\cal_pd270[1]~q ),
	.datae(!\cal_inc[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add9~0 .extended_lut = "off";
defparam \Add9~0 .lut_mask = 64'h3336933333369333;
defparam \Add9~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h0000FFFF00000000;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector34~0 (
	.dataa(!\cal_done[3]~q ),
	.datab(!\cal_pd270[3]~q ),
	.datac(!\cal_pd270~0_combout ),
	.datad(!\cal_pd270~2_combout ),
	.datae(!\Add9~0_combout ),
	.dataf(!\Add3~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector34~0 .extended_lut = "off";
defparam \Selector34~0 .lut_mask = 64'hCEF0C4F0CE00C400;
defparam \Selector34~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector34~1 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\cal_pd270[3]~q ),
	.datad(!\Selector34~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector34~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector34~1 .extended_lut = "off";
defparam \Selector34~1 .lut_mask = 64'h3B083B083B083B08;
defparam \Selector34~1 .shared_arith = "off";

dffeas \cal_pd270[3] (
	.clk(clock),
	.d(\Selector34~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_pd270[3]~q ),
	.prn(vcc));
defparam \cal_pd270[3] .is_wysiwyg = "true";
defparam \cal_pd270[3] .power_up = "low";

cyclonev_lcell_comb \Selector62~0 (
	.dataa(!\cal_pd270[3]~q ),
	.datab(!\cal_inc[3]~q ),
	.datac(!\cal_pd270_l[3]~q ),
	.datad(!\edges[3]~0_combout ),
	.datae(!\Equal10~0_combout ),
	.dataf(!\cal_pd270~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector62~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector62~0 .extended_lut = "off";
defparam \Selector62~0 .lut_mask = 64'h00FF00DE00000000;
defparam \Selector62~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector62~1 (
	.dataa(!\cal_done[3]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\WideOr8~0_combout ),
	.datad(!\Selector57~2_combout ),
	.datae(!\ignore_solid[3]~q ),
	.dataf(!\Selector62~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector62~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector62~1 .extended_lut = "off";
defparam \Selector62~1 .lut_mask = 64'hE000FFFFC000DDDD;
defparam \Selector62~1 .shared_arith = "off";

dffeas \ignore_solid[3] (
	.clk(clock),
	.d(\Selector62~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ignore_solid[3]~q ),
	.prn(vcc));
defparam \ignore_solid[3] .is_wysiwyg = "true";
defparam \ignore_solid[3] .power_up = "low";

dffeas \data_e0q[3] (
	.clk(clock),
	.d(\pd270_det|ff2~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e0q[3]~q ),
	.prn(vcc));
defparam \data_e0q[3] .is_wysiwyg = "true";
defparam \data_e0q[3] .power_up = "low";

dffeas \data_e1q[3] (
	.clk(clock),
	.d(\data_e0q[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\data_e1q[3]~q ),
	.prn(vcc));
defparam \data_e1q[3] .is_wysiwyg = "true";
defparam \data_e1q[3] .power_up = "low";

cyclonev_lcell_comb \edges[3]~0 (
	.dataa(!\pd_0_p[3]~q ),
	.datab(!\pd_0[3]~q ),
	.datac(!\pd_1_p[3]~q ),
	.datad(!\pd_1[3]~q ),
	.datae(!\ignore_solid[3]~q ),
	.dataf(!\data_e1q[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\edges[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \edges[3]~0 .extended_lut = "off";
defparam \edges[3]~0 .lut_mask = 64'hF99FFFFF00000000;
defparam \edges[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector54~0 (
	.dataa(!\cal_done[3]~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\Selector56~0_combout ),
	.datad(!\edges[3]~0_combout ),
	.datae(!\cal_pd270~0_combout ),
	.dataf(!\cal_pd270~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector54~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector54~0 .extended_lut = "off";
defparam \Selector54~0 .lut_mask = 64'h7373505073735073;
defparam \Selector54~0 .shared_arith = "off";

dffeas \cal_done[3] (
	.clk(clock),
	.d(\Selector54~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_done[3]~q ),
	.prn(vcc));
defparam \cal_done[3] .is_wysiwyg = "true";
defparam \cal_done[3] .power_up = "low";

cyclonev_lcell_comb WideAnd0(
	.dataa(!\cal_done[0]~q ),
	.datab(!\cal_done[1]~q ),
	.datac(!\cal_done[2]~q ),
	.datad(!\cal_done[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideAnd0.extended_lut = "off";
defparam WideAnd0.lut_mask = 64'h0001000100010001;
defparam WideAnd0.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\state.IDLE~q ),
	.datab(!\Equal11~2_combout ),
	.datac(!\state.TESTBUS_SET~q ),
	.datad(!\cal_en~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h0C530C530C530C53;
defparam \Selector0~0 .shared_arith = "off";

dffeas cal_en(
	.clk(clock),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\cal_en~q ),
	.prn(vcc));
defparam cal_en.is_wysiwyg = "true";
defparam cal_en.power_up = "low";

cyclonev_lcell_comb \Selector83~0 (
	.dataa(!\state.PDOF_TEST_WR~q ),
	.datab(!\ret_state.CAL_PD_WR~q ),
	.datac(!\Selector82~0_combout ),
	.datad(!\cal_en~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector83~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector83~0 .extended_lut = "off";
defparam \Selector83~0 .lut_mask = 64'h0357035703570357;
defparam \Selector83~0 .shared_arith = "off";

dffeas \ret_state.CAL_PD_WR (
	.clk(clock),
	.d(\Selector83~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ret_state.CAL_PD_WR~q ),
	.prn(vcc));
defparam \ret_state.CAL_PD_WR .is_wysiwyg = "true";
defparam \ret_state.CAL_PD_WR .power_up = "low";

cyclonev_lcell_comb \Selector14~0 (
	.dataa(!\state~25_combout ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\WideAnd0~combout ),
	.datad(!\ret_state.CAL_PD_WR~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~0 .extended_lut = "off";
defparam \Selector14~0 .lut_mask = 64'h3075307530753075;
defparam \Selector14~0 .shared_arith = "off";

dffeas \state.CAL_PD_WR (
	.clk(clock),
	.d(\Selector14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CAL_PD_WR~q ),
	.prn(vcc));
defparam \state.CAL_PD_WR .is_wysiwyg = "true";
defparam \state.CAL_PD_WR .power_up = "low";

cyclonev_lcell_comb \WideAnd1~0 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_done[0]~q ),
	.datac(!\cal_done[1]~q ),
	.datad(!\cal_done[2]~q ),
	.datae(!\cal_done[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideAnd1~0 .extended_lut = "off";
defparam \WideAnd1~0 .lut_mask = 64'h0000000100000001;
defparam \WideAnd1~0 .shared_arith = "off";

cyclonev_lcell_comb \WideAnd1~1 (
	.dataa(!\cal_pd0[0]~q ),
	.datab(!\cal_pd0[3]~q ),
	.datac(!\cal_pd0[2]~q ),
	.datad(!\cal_pd0[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideAnd1~1 .extended_lut = "off";
defparam \WideAnd1~1 .lut_mask = 64'h8001800180018001;
defparam \WideAnd1~1 .shared_arith = "off";

cyclonev_lcell_comb \WideAnd2~0 (
	.dataa(!\cal_pd180[3]~q ),
	.datab(!\cal_pd180[2]~q ),
	.datac(!\cal_pd180[1]~q ),
	.datad(!\cal_pd180[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideAnd2~0 .extended_lut = "off";
defparam \WideAnd2~0 .lut_mask = 64'h8001800180018001;
defparam \WideAnd2~0 .shared_arith = "off";

cyclonev_lcell_comb \WideAnd3~0 (
	.dataa(!\cal_pd270[0]~q ),
	.datab(!\cal_pd270[3]~q ),
	.datac(!\cal_pd270[2]~q ),
	.datad(!\cal_pd270[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideAnd3~0 .extended_lut = "off";
defparam \WideAnd3~0 .lut_mask = 64'h8001800180018001;
defparam \WideAnd3~0 .shared_arith = "off";

cyclonev_lcell_comb \WideAnd4~0 (
	.dataa(!\cal_pd90[3]~q ),
	.datab(!\cal_pd90[2]~q ),
	.datac(!\cal_pd90[1]~q ),
	.datad(!\cal_pd90[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideAnd4~0 .extended_lut = "off";
defparam \WideAnd4~0 .lut_mask = 64'h8001800180018001;
defparam \WideAnd4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~0 (
	.dataa(!\WideAnd1~1_combout ),
	.datab(!\WideAnd2~0_combout ),
	.datac(!\WideAnd3~0_combout ),
	.datad(!\WideAnd4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~0 .extended_lut = "off";
defparam \Selector75~0 .lut_mask = 64'h8000800080008000;
defparam \Selector75~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~1 (
	.dataa(!\state.SAMPLE_TB~q ),
	.datab(!\recal_counter[0]~q ),
	.datac(!\recal_counter[1]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~1 .extended_lut = "off";
defparam \Selector75~1 .lut_mask = 64'h5555550155555501;
defparam \Selector75~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~2 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\state.CH_WAIT~q ),
	.datac(!\WideAnd0~combout ),
	.datad(!\state.SAMPLE_TB~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~2 .extended_lut = "off";
defparam \Selector75~2 .lut_mask = 64'hD850D850D850D850;
defparam \Selector75~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector75~3 (
	.dataa(!\WideAnd1~0_combout ),
	.datab(!\do_recal~q ),
	.datac(!\Selector75~0_combout ),
	.datad(!\Selector75~1_combout ),
	.datae(!\Selector75~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~3 .extended_lut = "off";
defparam \Selector75~3 .lut_mask = 64'h5073737350737373;
defparam \Selector75~3 .shared_arith = "off";

dffeas do_recal(
	.clk(clock),
	.d(\Selector75~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\do_recal~q ),
	.prn(vcc));
defparam do_recal.is_wysiwyg = "true";
defparam do_recal.power_up = "low";

cyclonev_lcell_comb \always1~0 (
	.dataa(!\do_recal~q ),
	.datab(!\recal_counter[0]~q ),
	.datac(!\recal_counter[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'h5454545454545454;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \counter[2]~1 (
	.dataa(!reset),
	.datab(!\state.CH_WAIT~q ),
	.datac(!\state.SAMPLE_TB~q ),
	.datad(!\always1~0_combout ),
	.datae(!\Equal1~1_combout ),
	.dataf(!\state.DPRIO_WAIT~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter[2]~1 .extended_lut = "off";
defparam \counter[2]~1 .lut_mask = 64'hBFBFBABFFFFFFAFF;
defparam \counter[2]~1 .shared_arith = "off";

dffeas \counter[3] (
	.clk(clock),
	.d(\Add4~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[3]~q ),
	.prn(vcc));
defparam \counter[3] .is_wysiwyg = "true";
defparam \counter[3] .power_up = "low";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~13 .shared_arith = "off";

dffeas \counter[4] (
	.clk(clock),
	.d(\Add4~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[4]~q ),
	.prn(vcc));
defparam \counter[4] .is_wysiwyg = "true";
defparam \counter[4] .power_up = "low";

cyclonev_lcell_comb \Add4~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~29_sumout ),
	.cout(\Add4~30 ),
	.shareout());
defparam \Add4~29 .extended_lut = "off";
defparam \Add4~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~29 .shared_arith = "off";

dffeas \counter[5] (
	.clk(clock),
	.d(\Add4~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[5]~q ),
	.prn(vcc));
defparam \counter[5] .is_wysiwyg = "true";
defparam \counter[5] .power_up = "low";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~25_sumout ),
	.cout(\Add4~26 ),
	.shareout());
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~25 .shared_arith = "off";

dffeas \counter[6] (
	.clk(clock),
	.d(\Add4~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[6]~q ),
	.prn(vcc));
defparam \counter[6] .is_wysiwyg = "true";
defparam \counter[6] .power_up = "low";

cyclonev_lcell_comb \pd_0_p[0]~0 (
	.dataa(!\counter[1]~q ),
	.datab(!\counter[6]~q ),
	.datac(!\counter[5]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\state.DPRIO_WAIT~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_0_p[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_0_p[0]~0 .extended_lut = "off";
defparam \pd_0_p[0]~0 .lut_mask = 64'h0000004000000040;
defparam \pd_0_p[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \counter[2]~0 (
	.dataa(!reset),
	.datab(!\state.CH_WAIT~q ),
	.datac(!\state.SAMPLE_TB~q ),
	.datad(!\Equal1~1_combout ),
	.datae(!\pd_0_p[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter[2]~0 .extended_lut = "off";
defparam \counter[2]~0 .lut_mask = 64'hBBBFFFFFBBBFFFFF;
defparam \counter[2]~0 .shared_arith = "off";

dffeas \counter[0] (
	.clk(clock),
	.d(\Add4~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[0]~q ),
	.prn(vcc));
defparam \counter[0] .is_wysiwyg = "true";
defparam \counter[0] .power_up = "low";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(\Add4~22 ),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~21 .shared_arith = "off";

dffeas \counter[1] (
	.clk(clock),
	.d(\Add4~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[1]~q ),
	.prn(vcc));
defparam \counter[1] .is_wysiwyg = "true";
defparam \counter[1] .power_up = "low";

dffeas \counter[2] (
	.clk(clock),
	.d(\Add4~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[2]~q ),
	.prn(vcc));
defparam \counter[2] .is_wysiwyg = "true";
defparam \counter[2] .power_up = "low";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~9 .shared_arith = "off";

dffeas \counter[7] (
	.clk(clock),
	.d(\Add4~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter[2]~0_combout ),
	.sload(gnd),
	.ena(\counter[2]~1_combout ),
	.q(\counter[7]~q ),
	.prn(vcc));
defparam \counter[7] .is_wysiwyg = "true";
defparam \counter[7] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\counter[2]~q ),
	.datab(!\counter[0]~q ),
	.datac(!\counter[7]~q ),
	.datad(!\counter[4]~q ),
	.datae(!\counter[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h4000000040000000;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'h1111111111111111;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!\state.SAMPLE_TB~q ),
	.datab(!\Equal1~1_combout ),
	.datac(!\pd_0_p[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'h4F4F4F4F4F4F4F4F;
defparam \Selector16~0 .shared_arith = "off";

dffeas \state.SAMPLE_TB (
	.clk(clock),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.SAMPLE_TB~q ),
	.prn(vcc));
defparam \state.SAMPLE_TB .is_wysiwyg = "true";
defparam \state.SAMPLE_TB .power_up = "low";

cyclonev_lcell_comb \state~30 (
	.dataa(!reset),
	.datab(!\state.SAMPLE_TB~q ),
	.datac(!\Equal1~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~30 .extended_lut = "off";
defparam \state~30 .lut_mask = 64'h0101010101010101;
defparam \state~30 .shared_arith = "off";

dffeas \state.TEST_INPUT (
	.clk(clock),
	.d(\state~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.TEST_INPUT~q ),
	.prn(vcc));
defparam \state.TEST_INPUT .is_wysiwyg = "true";
defparam \state.TEST_INPUT .power_up = "low";

cyclonev_lcell_comb \Selector13~0 (
	.dataa(!\state.CH_WAIT~q ),
	.datab(!\state.TEST_INPUT~q ),
	.datac(!\WideAnd0~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~0 .extended_lut = "off";
defparam \Selector13~0 .lut_mask = 64'h5757575757575757;
defparam \Selector13~0 .shared_arith = "off";

dffeas \state.TESTBUS_SET (
	.clk(clock),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.TESTBUS_SET~q ),
	.prn(vcc));
defparam \state.TESTBUS_SET .is_wysiwyg = "true";
defparam \state.TESTBUS_SET .power_up = "low";

cyclonev_lcell_comb \state~29 (
	.dataa(!reset),
	.datab(!\Equal11~2_combout ),
	.datac(!\state.TESTBUS_SET~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~29 .extended_lut = "off";
defparam \state~29 .lut_mask = 64'h0404040404040404;
defparam \state~29 .shared_arith = "off";

dffeas \state.CHECK_PLL_RD (
	.clk(clock),
	.d(\state~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CHECK_PLL_RD~q ),
	.prn(vcc));
defparam \state.CHECK_PLL_RD .is_wysiwyg = "true";
defparam \state.CHECK_PLL_RD .power_up = "low";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!\state.CHECK_PLL_RD~q ),
	.datab(!\state.PDOF_TEST_RD~q ),
	.datac(!alt_cal_dprio_datain_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \Selector18~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~1 (
	.dataa(!read1),
	.datab(!\Equal11~2_combout ),
	.datac(!\state.DPRIO_READ~q ),
	.datad(!\state~28_combout ),
	.datae(!\Selector18~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~1 .extended_lut = "off";
defparam \Selector18~1 .lut_mask = 64'hFFFF0F04FFFF0F04;
defparam \Selector18~1 .shared_arith = "off";

dffeas \state.DPRIO_READ (
	.clk(clock),
	.d(\Selector18~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.DPRIO_READ~q ),
	.prn(vcc));
defparam \state.DPRIO_READ .is_wysiwyg = "true";
defparam \state.DPRIO_READ .power_up = "low";

cyclonev_lcell_comb \state~25 (
	.dataa(!write_reg1),
	.datab(!read1),
	.datac(!\state.DPRIO_WRITE~q ),
	.datad(!alt_cal_dprio_busy),
	.datae(!\did_dprio~q ),
	.dataf(!\state.DPRIO_READ~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~25 .extended_lut = "off";
defparam \state~25 .lut_mask = 64'h00000A000000CE00;
defparam \state~25 .shared_arith = "off";

cyclonev_lcell_comb \Selector87~0 (
	.dataa(!\state.PDOF_TEST_RD~q ),
	.datab(!\ret_state.PDOF_TEST_WR~q ),
	.datac(!\Selector82~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector87~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector87~0 .extended_lut = "off";
defparam \Selector87~0 .lut_mask = 64'h5757575757575757;
defparam \Selector87~0 .shared_arith = "off";

dffeas \ret_state.PDOF_TEST_WR (
	.clk(clock),
	.d(\Selector87~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ret_state.PDOF_TEST_WR~q ),
	.prn(vcc));
defparam \ret_state.PDOF_TEST_WR .is_wysiwyg = "true";
defparam \ret_state.PDOF_TEST_WR .power_up = "low";

cyclonev_lcell_comb \Selector21~0 (
	.dataa(!\state~25_combout ),
	.datab(!\ret_state.PDOF_TEST_WR~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~0 .extended_lut = "off";
defparam \Selector21~0 .lut_mask = 64'h1111111111111111;
defparam \Selector21~0 .shared_arith = "off";

dffeas \state.PDOF_TEST_WR (
	.clk(clock),
	.d(\Selector21~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.PDOF_TEST_WR~q ),
	.prn(vcc));
defparam \state.PDOF_TEST_WR .is_wysiwyg = "true";
defparam \state.PDOF_TEST_WR .power_up = "low";

cyclonev_lcell_comb \Selector104~0 (
	.dataa(!\state.PDOF_TEST_WR~q ),
	.datab(!\state.CAL_PD_WR~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector104~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector104~0 .extended_lut = "off";
defparam \Selector104~0 .lut_mask = 64'h8888888888888888;
defparam \Selector104~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!write_reg1),
	.datab(!\state.DPRIO_WRITE~q ),
	.datac(!\Selector104~0_combout ),
	.datad(!\Equal11~2_combout ),
	.datae(!\state~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'hF3F3F1F0F3F3F1F0;
defparam \Selector19~0 .shared_arith = "off";

dffeas \state.DPRIO_WRITE (
	.clk(clock),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.DPRIO_WRITE~q ),
	.prn(vcc));
defparam \state.DPRIO_WRITE .is_wysiwyg = "true";
defparam \state.DPRIO_WRITE .power_up = "low";

cyclonev_lcell_comb \Selector82~1 (
	.dataa(!\state.DPRIO_WRITE~q ),
	.datab(!alt_cal_dprio_busy),
	.datac(!\did_dprio~q ),
	.datad(!\state.DPRIO_READ~q ),
	.datae(!\Selector82~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector82~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector82~1 .extended_lut = "off";
defparam \Selector82~1 .lut_mask = 64'h45CF4FCF45CF4FCF;
defparam \Selector82~1 .shared_arith = "off";

dffeas did_dprio(
	.clk(clock),
	.d(\Selector82~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\did_dprio~q ),
	.prn(vcc));
defparam did_dprio.is_wysiwyg = "true";
defparam did_dprio.power_up = "low";

cyclonev_lcell_comb \state~28 (
	.dataa(!alt_cal_dprio_busy),
	.datab(!\did_dprio~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~28 .extended_lut = "off";
defparam \state~28 .lut_mask = 64'h2222222222222222;
defparam \state~28 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!\state.PDOF_TEST_RD~q ),
	.datab(!alt_cal_dprio_datain_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'h1111111111111111;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~1 (
	.dataa(!write_reg1),
	.datab(!read1),
	.datac(!\state.DPRIO_WRITE~q ),
	.datad(!\state.DPRIO_READ~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~1 .extended_lut = "off";
defparam \Selector17~1 .lut_mask = 64'h0537053705370537;
defparam \Selector17~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector85~0 (
	.dataa(!\state.PDOF_TEST_WR~q ),
	.datab(!\Selector82~0_combout ),
	.datac(!\ret_state.CH_ADV~q ),
	.datad(!\cal_en~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector85~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector85~0 .extended_lut = "off";
defparam \Selector85~0 .lut_mask = 64'h5703570357035703;
defparam \Selector85~0 .shared_arith = "off";

dffeas \ret_state.CH_ADV (
	.clk(clock),
	.d(\Selector85~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\ret_state.CH_ADV~q ),
	.prn(vcc));
defparam \ret_state.CH_ADV .is_wysiwyg = "true";
defparam \ret_state.CH_ADV .power_up = "low";

cyclonev_lcell_comb \Selector17~2 (
	.dataa(!write_reg1),
	.datab(!read1),
	.datac(!\state.DPRIO_WRITE~q ),
	.datad(!\state.DPRIO_READ~q ),
	.datae(!\ret_state.CH_ADV~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~2 .extended_lut = "off";
defparam \Selector17~2 .lut_mask = 64'h00000ACE00000ACE;
defparam \Selector17~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~3 (
	.dataa(!\Equal11~2_combout ),
	.datab(!\state~28_combout ),
	.datac(!\state.TESTBUS_SET~q ),
	.datad(!\Selector17~0_combout ),
	.datae(!\Selector17~1_combout ),
	.dataf(!\Selector17~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~3 .extended_lut = "off";
defparam \Selector17~3 .lut_mask = 64'h05FF15FF37FF37FF;
defparam \Selector17~3 .shared_arith = "off";

dffeas \state.CH_ADV (
	.clk(clock),
	.d(\Selector17~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\state.CH_ADV~q ),
	.prn(vcc));
defparam \state.CH_ADV .is_wysiwyg = "true";
defparam \state.CH_ADV .power_up = "low";

cyclonev_lcell_comb \ret_state~12 (
	.dataa(!reset),
	.datab(!\ret_state.IDLE~q ),
	.datac(!\Selector82~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ret_state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ret_state~12 .extended_lut = "off";
defparam \ret_state~12 .lut_mask = 64'h5151515151515151;
defparam \ret_state~12 .shared_arith = "off";

dffeas \ret_state.IDLE (
	.clk(clock),
	.d(\ret_state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ret_state.IDLE~q ),
	.prn(vcc));
defparam \ret_state.IDLE .is_wysiwyg = "true";
defparam \ret_state.IDLE .power_up = "low";

cyclonev_lcell_comb \state~26 (
	.dataa(!reset),
	.datab(!\state.IDLE~q ),
	.datac(!\Selector11~0_combout ),
	.datad(!\ret_state.IDLE~q ),
	.datae(!\state~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~26 .extended_lut = "off";
defparam \state~26 .lut_mask = 64'h1515001515150015;
defparam \state~26 .shared_arith = "off";

cyclonev_lcell_comb \state~27 (
	.dataa(!alt_cal_channel_9),
	.datab(!\LessThan1~2_combout ),
	.datac(!\state.CH_ADV~q ),
	.datad(!\state~26_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~27 .extended_lut = "off";
defparam \state~27 .lut_mask = 64'h00F200F200F200F2;
defparam \state~27 .shared_arith = "off";

dffeas \state.IDLE (
	.clk(clock),
	.d(\state~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.IDLE~q ),
	.prn(vcc));
defparam \state.IDLE .is_wysiwyg = "true";
defparam \state.IDLE .power_up = "low";

cyclonev_lcell_comb \alt_cal_busy~0 (
	.dataa(!alt_cal_busy1),
	.datab(!\state.IDLE~q ),
	.datac(!\Selector11~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\alt_cal_busy~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \alt_cal_busy~0 .extended_lut = "off";
defparam \alt_cal_busy~0 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \alt_cal_busy~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector104~1 (
	.dataa(!write_reg1),
	.datab(!\state.DPRIO_WRITE~q ),
	.datac(!\Selector104~0_combout ),
	.datad(!alt_cal_dprio_busy),
	.datae(!\did_dprio~q ),
	.dataf(!\Equal11~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector104~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector104~1 .extended_lut = "off";
defparam \Selector104~1 .lut_mask = 64'h3704150437040404;
defparam \Selector104~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector81~1 (
	.dataa(!read1),
	.datab(!alt_cal_dprio_busy),
	.datac(!\did_dprio~q ),
	.datad(!\Equal11~2_combout ),
	.datae(!\state.DPRIO_READ~q ),
	.dataf(!\Selector81~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector81~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector81~1 .extended_lut = "off";
defparam \Selector81~1 .lut_mask = 64'h0000C4C05555C4C0;
defparam \Selector81~1 .shared_arith = "off";

cyclonev_lcell_comb \Add10~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~17_sumout ),
	.cout(\Add10~18 ),
	.shareout());
defparam \Add10~17 .extended_lut = "off";
defparam \Add10~17 .lut_mask = 64'h00000000000000FF;
defparam \Add10~17 .shared_arith = "off";

cyclonev_lcell_comb \Add10~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~21_sumout ),
	.cout(\Add10~22 ),
	.shareout());
defparam \Add10~21 .extended_lut = "off";
defparam \Add10~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~21 .shared_arith = "off";

cyclonev_lcell_comb \Add10~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~25_sumout ),
	.cout(\Add10~26 ),
	.shareout());
defparam \Add10~25 .extended_lut = "off";
defparam \Add10~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~25 .shared_arith = "off";

cyclonev_lcell_comb \Add10~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~29_sumout ),
	.cout(\Add10~30 ),
	.shareout());
defparam \Add10~29 .extended_lut = "off";
defparam \Add10~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~29 .shared_arith = "off";

cyclonev_lcell_comb \Add10~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~33_sumout ),
	.cout(\Add10~34 ),
	.shareout());
defparam \Add10~33 .extended_lut = "off";
defparam \Add10~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~33 .shared_arith = "off";

cyclonev_lcell_comb \Add10~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~37_sumout ),
	.cout(\Add10~38 ),
	.shareout());
defparam \Add10~37 .extended_lut = "off";
defparam \Add10~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~37 .shared_arith = "off";

cyclonev_lcell_comb \Add10~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~5_sumout ),
	.cout(\Add10~6 ),
	.shareout());
defparam \Add10~5 .extended_lut = "off";
defparam \Add10~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~5 .shared_arith = "off";

cyclonev_lcell_comb \Add10~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~9_sumout ),
	.cout(\Add10~10 ),
	.shareout());
defparam \Add10~9 .extended_lut = "off";
defparam \Add10~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~9 .shared_arith = "off";

cyclonev_lcell_comb \Add10~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~13_sumout ),
	.cout(\Add10~14 ),
	.shareout());
defparam \Add10~13 .extended_lut = "off";
defparam \Add10~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~13 .shared_arith = "off";

cyclonev_lcell_comb \Add10~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!alt_cal_channel_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~1_sumout ),
	.cout(),
	.shareout());
defparam \Add10~1 .extended_lut = "off";
defparam \Add10~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add10~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!alt_cal_channel_9),
	.datab(!\state.IDLE~q ),
	.datac(!\LessThan1~2_combout ),
	.datad(!\state.CH_ADV~q ),
	.datae(!\Add10~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h1155115F1155115F;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!\state.IDLE~q ),
	.datab(!\state.CH_ADV~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h8888888888888888;
defparam \Selector10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!alt_cal_channel_6),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~5_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h5073507350735073;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!alt_cal_channel_7),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~9_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h5073507350735073;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!alt_cal_channel_8),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~13_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h5073507350735073;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~1 (
	.dataa(!alt_cal_channel_0),
	.datab(!\Add10~17_sumout ),
	.datac(!\Selector12~0_combout ),
	.datad(!\Selector10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~1 .extended_lut = "off";
defparam \Selector10~1 .lut_mask = 64'h5703570357035703;
defparam \Selector10~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!alt_cal_channel_1),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~21_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h5073507350735073;
defparam \Selector9~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!alt_cal_channel_2),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h5073507350735073;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!alt_cal_channel_3),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~29_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h5073507350735073;
defparam \Selector7~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!alt_cal_channel_4),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~33_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h5073507350735073;
defparam \Selector6~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!alt_cal_channel_5),
	.datab(!\Selector12~0_combout ),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add10~37_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h5073507350735073;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector79~0 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\Selector81~0_combout ),
	.datac(!address_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector79~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector79~0 .extended_lut = "off";
defparam \Selector79~0 .lut_mask = 64'h5757575757575757;
defparam \Selector79~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector80~0 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\state.CHECK_PLL_RD~q ),
	.datac(!\state.PDOF_TEST_RD~q ),
	.datad(!address_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector80~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector80~0 .extended_lut = "off";
defparam \Selector80~0 .lut_mask = 64'h77F777F777F777F7;
defparam \Selector80~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector76~0 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\Selector81~0_combout ),
	.datac(!address_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~0 .extended_lut = "off";
defparam \Selector76~0 .lut_mask = 64'hCECECECECECECECE;
defparam \Selector76~0 .shared_arith = "off";

cyclonev_lcell_comb \dataout[0]~0 (
	.dataa(!reset),
	.datab(!\WideAnd1~0_combout ),
	.datac(!\WideAnd1~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout[0]~0 .extended_lut = "off";
defparam \dataout[0]~0 .lut_mask = 64'h5454545454545454;
defparam \dataout[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dataout~1 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd0[3]~q ),
	.datac(!\cal_pd0[1]~q ),
	.datad(!\dataout[0]~0_combout ),
	.datae(!alt_cal_dprio_datain_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~1 .extended_lut = "off";
defparam \dataout~1 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~1 .shared_arith = "off";

cyclonev_lcell_comb \dataout[0]~2 (
	.dataa(!reset),
	.datab(!\state.PDOF_TEST_WR~q ),
	.datac(!\state.CAL_PD_WR~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout[0]~2 .extended_lut = "off";
defparam \dataout[0]~2 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \dataout[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \dataout~3 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd0[3]~q ),
	.datac(!\cal_pd0[2]~q ),
	.datad(!\dataout[0]~0_combout ),
	.datae(!\cal_en~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~3 .extended_lut = "off";
defparam \dataout~3 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~3 .shared_arith = "off";

cyclonev_lcell_comb \dataout~4 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd0[0]~q ),
	.datac(!\cal_pd0[3]~q ),
	.datad(!\dataout[0]~0_combout ),
	.datae(!alt_cal_dprio_datain_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~4 .extended_lut = "off";
defparam \dataout~4 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~4 .shared_arith = "off";

cyclonev_lcell_comb \dataout~5 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd0[3]~q ),
	.datac(!\dataout[0]~0_combout ),
	.datad(!alt_cal_dprio_datain_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~5 .extended_lut = "off";
defparam \dataout~5 .lut_mask = 64'h040E040E040E040E;
defparam \dataout~5 .shared_arith = "off";

cyclonev_lcell_comb \dataout[5]~6 (
	.dataa(!reset),
	.datab(!\WideAnd1~0_combout ),
	.datac(!\WideAnd2~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout[5]~6 .extended_lut = "off";
defparam \dataout[5]~6 .lut_mask = 64'h5454545454545454;
defparam \dataout[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \dataout~7 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd180[3]~q ),
	.datac(!\cal_pd180[0]~q ),
	.datad(!\dataout[5]~6_combout ),
	.datae(!alt_cal_dprio_datain_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~7 .extended_lut = "off";
defparam \dataout~7 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~7 .shared_arith = "off";

cyclonev_lcell_comb \dataout~8 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd180[3]~q ),
	.datac(!\cal_pd180[1]~q ),
	.datad(!\dataout[5]~6_combout ),
	.datae(!alt_cal_dprio_datain_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~8 .extended_lut = "off";
defparam \dataout~8 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~8 .shared_arith = "off";

cyclonev_lcell_comb \dataout~9 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd180[3]~q ),
	.datac(!\cal_pd180[2]~q ),
	.datad(!\dataout[5]~6_combout ),
	.datae(!alt_cal_dprio_datain_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~9 .extended_lut = "off";
defparam \dataout~9 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~9 .shared_arith = "off";

cyclonev_lcell_comb \dataout~10 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd180[3]~q ),
	.datac(!\dataout[5]~6_combout ),
	.datad(!alt_cal_dprio_datain_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~10 .extended_lut = "off";
defparam \dataout~10 .lut_mask = 64'h040E040E040E040E;
defparam \dataout~10 .shared_arith = "off";

cyclonev_lcell_comb \dataout[8]~11 (
	.dataa(!reset),
	.datab(!\WideAnd1~0_combout ),
	.datac(!\WideAnd3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout[8]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout[8]~11 .extended_lut = "off";
defparam \dataout[8]~11 .lut_mask = 64'h5454545454545454;
defparam \dataout[8]~11 .shared_arith = "off";

cyclonev_lcell_comb \dataout~12 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd270[0]~q ),
	.datac(!\cal_pd270[3]~q ),
	.datad(!\dataout[8]~11_combout ),
	.datae(!alt_cal_dprio_datain_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~12 .extended_lut = "off";
defparam \dataout~12 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~12 .shared_arith = "off";

cyclonev_lcell_comb \dataout~13 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd270[3]~q ),
	.datac(!\cal_pd270[1]~q ),
	.datad(!\dataout[8]~11_combout ),
	.datae(!alt_cal_dprio_datain_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~13 .extended_lut = "off";
defparam \dataout~13 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~13 .shared_arith = "off";

cyclonev_lcell_comb \dataout~14 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd270[3]~q ),
	.datac(!\cal_pd270[2]~q ),
	.datad(!\dataout[8]~11_combout ),
	.datae(!alt_cal_dprio_datain_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~14 .extended_lut = "off";
defparam \dataout~14 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~14 .shared_arith = "off";

cyclonev_lcell_comb \dataout~15 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd270[3]~q ),
	.datac(!\dataout[8]~11_combout ),
	.datad(!alt_cal_dprio_datain_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~15 .extended_lut = "off";
defparam \dataout~15 .lut_mask = 64'h040E040E040E040E;
defparam \dataout~15 .shared_arith = "off";

cyclonev_lcell_comb \dataout[13]~16 (
	.dataa(!reset),
	.datab(!\WideAnd1~0_combout ),
	.datac(!\WideAnd4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout[13]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout[13]~16 .extended_lut = "off";
defparam \dataout[13]~16 .lut_mask = 64'h5454545454545454;
defparam \dataout[13]~16 .shared_arith = "off";

cyclonev_lcell_comb \dataout~17 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd90[3]~q ),
	.datac(!\cal_pd90[0]~q ),
	.datad(!\dataout[13]~16_combout ),
	.datae(!alt_cal_dprio_datain_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~17 .extended_lut = "off";
defparam \dataout~17 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~17 .shared_arith = "off";

cyclonev_lcell_comb \dataout~18 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd90[3]~q ),
	.datac(!\cal_pd90[1]~q ),
	.datad(!\dataout[13]~16_combout ),
	.datae(!alt_cal_dprio_datain_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~18 .extended_lut = "off";
defparam \dataout~18 .lut_mask = 64'h004100EB004100EB;
defparam \dataout~18 .shared_arith = "off";

cyclonev_lcell_comb \dataout~19 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!alt_cal_dprio_datain_14),
	.datac(!\cal_pd90[3]~q ),
	.datad(!\cal_pd90[2]~q ),
	.datae(!\dataout[13]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~19 .extended_lut = "off";
defparam \dataout~19 .lut_mask = 64'h0000722700007227;
defparam \dataout~19 .shared_arith = "off";

cyclonev_lcell_comb \dataout~20 (
	.dataa(!\state.CAL_PD_WR~q ),
	.datab(!\cal_pd90[3]~q ),
	.datac(!\dataout[13]~16_combout ),
	.datad(!alt_cal_dprio_datain_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dataout~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dataout~20 .extended_lut = "off";
defparam \dataout~20 .lut_mask = 64'h040E040E040E040E;
defparam \dataout~20 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_cal_edge_detect (
	reset,
	ff21,
	testbus)/* synthesis synthesis_greybox=0 */;
input 	reset;
output 	ff21;
input 	testbus;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_edge_det_ff1~q ;
wire \pd_xor~0_combout ;


dffeas ff2(
	.clk(\pd_xor~0_combout ),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ff21),
	.prn(vcc));
defparam ff2.is_wysiwyg = "true";
defparam ff2.power_up = "low";

dffeas alt_edge_det_ff1(
	.clk(!testbus),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\alt_edge_det_ff1~q ),
	.prn(vcc));
defparam alt_edge_det_ff1.is_wysiwyg = "true";
defparam alt_edge_det_ff1.power_up = "low";

cyclonev_lcell_comb \pd_xor~0 (
	.dataa(!\alt_edge_det_ff1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_xor~0 .extended_lut = "off";
defparam \pd_xor~0 .lut_mask = 64'h5555555555555555;
defparam \pd_xor~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_cal_edge_detect_1 (
	reset,
	ff21,
	testbus)/* synthesis synthesis_greybox=0 */;
input 	reset;
output 	ff21;
input 	testbus;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_edge_det_ff1~q ;
wire \pd_xor~0_combout ;


dffeas ff2(
	.clk(\pd_xor~0_combout ),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ff21),
	.prn(vcc));
defparam ff2.is_wysiwyg = "true";
defparam ff2.power_up = "low";

dffeas alt_edge_det_ff1(
	.clk(!testbus),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\alt_edge_det_ff1~q ),
	.prn(vcc));
defparam alt_edge_det_ff1.is_wysiwyg = "true";
defparam alt_edge_det_ff1.power_up = "low";

cyclonev_lcell_comb \pd_xor~0 (
	.dataa(!\alt_edge_det_ff1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_xor~0 .extended_lut = "off";
defparam \pd_xor~0 .lut_mask = 64'h5555555555555555;
defparam \pd_xor~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_cal_edge_detect_2 (
	reset,
	ff21,
	testbus)/* synthesis synthesis_greybox=0 */;
input 	reset;
output 	ff21;
input 	testbus;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_edge_det_ff1~q ;
wire \pd_xor~0_combout ;


dffeas ff2(
	.clk(\pd_xor~0_combout ),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ff21),
	.prn(vcc));
defparam ff2.is_wysiwyg = "true";
defparam ff2.power_up = "low";

dffeas alt_edge_det_ff1(
	.clk(!testbus),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\alt_edge_det_ff1~q ),
	.prn(vcc));
defparam alt_edge_det_ff1.is_wysiwyg = "true";
defparam alt_edge_det_ff1.power_up = "low";

cyclonev_lcell_comb \pd_xor~0 (
	.dataa(!\alt_edge_det_ff1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_xor~0 .extended_lut = "off";
defparam \pd_xor~0 .lut_mask = 64'h5555555555555555;
defparam \pd_xor~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_cal_edge_detect_3 (
	reset,
	ff21,
	testbus)/* synthesis synthesis_greybox=0 */;
input 	reset;
output 	ff21;
input 	testbus;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_edge_det_ff1~q ;
wire \pd_xor~0_combout ;


dffeas ff2(
	.clk(\pd_xor~0_combout ),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ff21),
	.prn(vcc));
defparam ff2.is_wysiwyg = "true";
defparam ff2.power_up = "low";

dffeas alt_edge_det_ff1(
	.clk(!testbus),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\alt_edge_det_ff1~q ),
	.prn(vcc));
defparam alt_edge_det_ff1.is_wysiwyg = "true";
defparam alt_edge_det_ff1.power_up = "low";

cyclonev_lcell_comb \pd_xor~0 (
	.dataa(!\alt_edge_det_ff1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pd_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pd_xor~0 .extended_lut = "off";
defparam \pd_xor~0 .lut_mask = 64'h5555555555555555;
defparam \pd_xor~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_altera_wait_generate_2 (
	resync_chains0sync_r_1,
	launch_reg1,
	wait_reg1,
	ifsel_notdone_resync,
	launch_signal,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
output 	launch_reg1;
output 	wait_reg1;
input 	ifsel_notdone_resync;
input 	launch_signal;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_reg~0_combout ;


RECONFIGURE_IP_alt_xcvr_resync_2 rst_sync(
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.clk(mgmt_clk_clk));

dffeas launch_reg(
	.clk(mgmt_clk_clk),
	.d(launch_signal),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(launch_reg1),
	.prn(vcc));
defparam launch_reg.is_wysiwyg = "true";
defparam launch_reg.power_up = "low";

dffeas wait_reg(
	.clk(mgmt_clk_clk),
	.d(\wait_reg~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_reg1),
	.prn(vcc));
defparam wait_reg.is_wysiwyg = "true";
defparam wait_reg.power_up = "low";

cyclonev_lcell_comb \wait_reg~0 (
	.dataa(!resync_chains0sync_r_1),
	.datab(!launch_signal),
	.datac(!launch_reg1),
	.datad(!wait_reg1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_reg~0 .extended_lut = "off";
defparam \wait_reg~0 .lut_mask = 64'h0100010001000100;
defparam \wait_reg~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_resync_2 (
	resync_chains0sync_r_1,
	ifsel_notdone_resync,
	clk)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
input 	ifsel_notdone_resync;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \resync_chains[0].sync_r[0]~q ;


dffeas \resync_chains[0].sync_r[1] (
	.clk(clk),
	.d(\resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resync_chains0sync_r_1),
	.prn(vcc));
defparam \resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[1] .power_up = "low";

dffeas \resync_chains[0].sync_r[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[0] .power_up = "low";

endmodule

module RECONFIGURE_IP_alt_xcvr_reconfig_pll (
	user_reconfig_readdata_10,
	user_reconfig_readdata_11,
	user_reconfig_readdata_12,
	basic_reconfig_readdata_12,
	user_reconfig_readdata_13,
	basic_reconfig_readdata_13,
	user_reconfig_readdata_14,
	basic_reconfig_readdata_14,
	user_reconfig_readdata_15,
	basic_reconfig_readdata_15,
	user_reconfig_readdata_16,
	basic_reconfig_readdata_16,
	user_reconfig_readdata_17,
	basic_reconfig_readdata_17,
	user_reconfig_readdata_18,
	basic_reconfig_readdata_18,
	user_reconfig_readdata_19,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	user_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	user_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	user_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	user_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	user_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	user_reconfig_readdata_0,
	Equal4,
	basic_reconfig_readdata_0,
	user_reconfig_readdata_1,
	basic_reconfig_readdata_1,
	user_reconfig_readdata_2,
	basic_reconfig_readdata_2,
	user_reconfig_readdata_3,
	basic_reconfig_readdata_3,
	user_reconfig_readdata_4,
	basic_reconfig_readdata_4,
	user_reconfig_readdata_5,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	user_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	user_reconfig_readdata_7,
	user_reconfig_readdata_8,
	basic_reconfig_readdata_8,
	user_reconfig_readdata_9,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	user_reconfig_readdata_25,
	user_reconfig_readdata_26,
	user_reconfig_readdata_27,
	user_reconfig_readdata_28,
	user_reconfig_readdata_29,
	user_reconfig_readdata_30,
	user_reconfig_readdata_31,
	master_write,
	grant_8,
	mutex_req,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	pll_mif_busy,
	ifsel_notdone_resync,
	uif_logical_ch_addr_0,
	comb,
	uif_logical_ch_addr_1,
	uif_logical_ch_addr_2,
	uif_logical_ch_addr_3,
	user_reconfig_readdata_101,
	uif_logical_ch_addr_4,
	uif_logical_ch_addr_5,
	uif_logical_ch_addr_6,
	uif_logical_ch_addr_7,
	uif_logical_ch_addr_8,
	uif_logical_ch_addr_9,
	mutex_grant,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	pll_go,
	uif_mode_0,
	Mux0,
	Mux3,
	WideOr0,
	pll_type,
	mif_rec_addr_7,
	mif_rec_addr_5,
	mif_rec_addr_6,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_10;
output 	user_reconfig_readdata_11;
output 	user_reconfig_readdata_12;
input 	basic_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
input 	basic_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
input 	basic_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
input 	basic_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
input 	basic_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
input 	basic_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
input 	basic_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
output 	user_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
output 	user_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
output 	user_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
output 	user_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
output 	user_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	user_reconfig_readdata_0;
input 	Equal4;
input 	basic_reconfig_readdata_0;
output 	user_reconfig_readdata_1;
input 	basic_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
input 	basic_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
input 	basic_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
input 	basic_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
output 	user_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
output 	user_reconfig_readdata_7;
output 	user_reconfig_readdata_8;
input 	basic_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	user_reconfig_readdata_25;
output 	user_reconfig_readdata_26;
output 	user_reconfig_readdata_27;
output 	user_reconfig_readdata_28;
output 	user_reconfig_readdata_29;
output 	user_reconfig_readdata_30;
output 	user_reconfig_readdata_31;
output 	master_write;
input 	grant_8;
output 	mutex_req;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
output 	pll_mif_busy;
input 	ifsel_notdone_resync;
input 	uif_logical_ch_addr_0;
input 	comb;
input 	uif_logical_ch_addr_1;
input 	uif_logical_ch_addr_2;
input 	uif_logical_ch_addr_3;
output 	user_reconfig_readdata_101;
input 	uif_logical_ch_addr_4;
input 	uif_logical_ch_addr_5;
input 	uif_logical_ch_addr_6;
input 	uif_logical_ch_addr_7;
input 	uif_logical_ch_addr_8;
input 	uif_logical_ch_addr_9;
output 	mutex_grant;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
output 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
input 	pll_go;
input 	uif_mode_0;
output 	Mux0;
output 	Mux3;
input 	WideOr0;
input 	pll_type;
input 	mif_rec_addr_7;
input 	mif_rec_addr_5;
input 	mif_rec_addr_6;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



RECONFIGURE_IP_av_xcvr_reconfig_pll pll_reconfig_av(
	.user_reconfig_readdata_10(user_reconfig_readdata_10),
	.user_reconfig_readdata_11(user_reconfig_readdata_11),
	.user_reconfig_readdata_12(user_reconfig_readdata_12),
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.user_reconfig_readdata_13(user_reconfig_readdata_13),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.user_reconfig_readdata_14(user_reconfig_readdata_14),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.user_reconfig_readdata_15(user_reconfig_readdata_15),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.user_reconfig_readdata_16(user_reconfig_readdata_16),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.user_reconfig_readdata_17(user_reconfig_readdata_17),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.user_reconfig_readdata_18(user_reconfig_readdata_18),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.user_reconfig_readdata_19(user_reconfig_readdata_19),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.user_reconfig_readdata_20(user_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.user_reconfig_readdata_21(user_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.user_reconfig_readdata_22(user_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.user_reconfig_readdata_23(user_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.user_reconfig_readdata_24(user_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.user_reconfig_readdata_0(user_reconfig_readdata_0),
	.Equal4(Equal4),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.user_reconfig_readdata_1(user_reconfig_readdata_1),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.user_reconfig_readdata_2(user_reconfig_readdata_2),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.user_reconfig_readdata_3(user_reconfig_readdata_3),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.user_reconfig_readdata_4(user_reconfig_readdata_4),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.user_reconfig_readdata_5(user_reconfig_readdata_5),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.user_reconfig_readdata_6(user_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.user_reconfig_readdata_7(user_reconfig_readdata_7),
	.user_reconfig_readdata_8(user_reconfig_readdata_8),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.user_reconfig_readdata_9(user_reconfig_readdata_9),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.user_reconfig_readdata_25(user_reconfig_readdata_25),
	.user_reconfig_readdata_26(user_reconfig_readdata_26),
	.user_reconfig_readdata_27(user_reconfig_readdata_27),
	.user_reconfig_readdata_28(user_reconfig_readdata_28),
	.user_reconfig_readdata_29(user_reconfig_readdata_29),
	.user_reconfig_readdata_30(user_reconfig_readdata_30),
	.user_reconfig_readdata_31(user_reconfig_readdata_31),
	.master_write(master_write),
	.grant_8(grant_8),
	.mutex_req(mutex_req),
	.master_address_2(master_address_2),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg(launch_reg),
	.wait_reg(wait_reg),
	.pll_mif_busy(pll_mif_busy),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.uif_logical_ch_addr_0(uif_logical_ch_addr_0),
	.comb(comb),
	.uif_logical_ch_addr_1(uif_logical_ch_addr_1),
	.uif_logical_ch_addr_2(uif_logical_ch_addr_2),
	.uif_logical_ch_addr_3(uif_logical_ch_addr_3),
	.user_reconfig_readdata_101(user_reconfig_readdata_101),
	.uif_logical_ch_addr_4(uif_logical_ch_addr_4),
	.uif_logical_ch_addr_5(uif_logical_ch_addr_5),
	.uif_logical_ch_addr_6(uif_logical_ch_addr_6),
	.uif_logical_ch_addr_7(uif_logical_ch_addr_7),
	.uif_logical_ch_addr_8(uif_logical_ch_addr_8),
	.uif_logical_ch_addr_9(uif_logical_ch_addr_9),
	.mutex_grant(mutex_grant),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.master_writedata_11(master_writedata_11),
	.master_writedata_12(master_writedata_12),
	.master_writedata_13(master_writedata_13),
	.master_writedata_14(master_writedata_14),
	.master_writedata_15(master_writedata_15),
	.pll_go(pll_go),
	.uif_mode_0(uif_mode_0),
	.Mux0(Mux0),
	.Mux3(Mux3),
	.WideOr0(WideOr0),
	.pll_type(pll_type),
	.mif_rec_addr_7(mif_rec_addr_7),
	.mif_rec_addr_5(mif_rec_addr_5),
	.mif_rec_addr_6(mif_rec_addr_6),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15));

endmodule

module RECONFIGURE_IP_av_xcvr_reconfig_pll (
	user_reconfig_readdata_10,
	user_reconfig_readdata_11,
	user_reconfig_readdata_12,
	basic_reconfig_readdata_12,
	user_reconfig_readdata_13,
	basic_reconfig_readdata_13,
	user_reconfig_readdata_14,
	basic_reconfig_readdata_14,
	user_reconfig_readdata_15,
	basic_reconfig_readdata_15,
	user_reconfig_readdata_16,
	basic_reconfig_readdata_16,
	user_reconfig_readdata_17,
	basic_reconfig_readdata_17,
	user_reconfig_readdata_18,
	basic_reconfig_readdata_18,
	user_reconfig_readdata_19,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	user_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	user_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	user_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	user_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	user_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	user_reconfig_readdata_0,
	Equal4,
	basic_reconfig_readdata_0,
	user_reconfig_readdata_1,
	basic_reconfig_readdata_1,
	user_reconfig_readdata_2,
	basic_reconfig_readdata_2,
	user_reconfig_readdata_3,
	basic_reconfig_readdata_3,
	user_reconfig_readdata_4,
	basic_reconfig_readdata_4,
	user_reconfig_readdata_5,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	user_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	user_reconfig_readdata_7,
	user_reconfig_readdata_8,
	basic_reconfig_readdata_8,
	user_reconfig_readdata_9,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	user_reconfig_readdata_25,
	user_reconfig_readdata_26,
	user_reconfig_readdata_27,
	user_reconfig_readdata_28,
	user_reconfig_readdata_29,
	user_reconfig_readdata_30,
	user_reconfig_readdata_31,
	master_write,
	grant_8,
	mutex_req,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	pll_mif_busy,
	ifsel_notdone_resync,
	uif_logical_ch_addr_0,
	comb,
	uif_logical_ch_addr_1,
	uif_logical_ch_addr_2,
	uif_logical_ch_addr_3,
	user_reconfig_readdata_101,
	uif_logical_ch_addr_4,
	uif_logical_ch_addr_5,
	uif_logical_ch_addr_6,
	uif_logical_ch_addr_7,
	uif_logical_ch_addr_8,
	uif_logical_ch_addr_9,
	mutex_grant,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	pll_go,
	uif_mode_0,
	Mux0,
	Mux3,
	WideOr0,
	pll_type,
	mif_rec_addr_7,
	mif_rec_addr_5,
	mif_rec_addr_6,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_10;
output 	user_reconfig_readdata_11;
output 	user_reconfig_readdata_12;
input 	basic_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
input 	basic_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
input 	basic_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
input 	basic_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
input 	basic_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
input 	basic_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
input 	basic_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
output 	user_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
output 	user_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
output 	user_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
output 	user_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
output 	user_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
output 	user_reconfig_readdata_0;
input 	Equal4;
input 	basic_reconfig_readdata_0;
output 	user_reconfig_readdata_1;
input 	basic_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
input 	basic_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
input 	basic_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
input 	basic_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
output 	user_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
output 	user_reconfig_readdata_7;
output 	user_reconfig_readdata_8;
input 	basic_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	user_reconfig_readdata_25;
output 	user_reconfig_readdata_26;
output 	user_reconfig_readdata_27;
output 	user_reconfig_readdata_28;
output 	user_reconfig_readdata_29;
output 	user_reconfig_readdata_30;
output 	user_reconfig_readdata_31;
output 	master_write;
input 	grant_8;
output 	mutex_req;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
output 	pll_mif_busy;
input 	ifsel_notdone_resync;
input 	uif_logical_ch_addr_0;
input 	comb;
input 	uif_logical_ch_addr_1;
input 	uif_logical_ch_addr_2;
input 	uif_logical_ch_addr_3;
output 	user_reconfig_readdata_101;
input 	uif_logical_ch_addr_4;
input 	uif_logical_ch_addr_5;
input 	uif_logical_ch_addr_6;
input 	uif_logical_ch_addr_7;
input 	uif_logical_ch_addr_8;
input 	uif_logical_ch_addr_9;
output 	mutex_grant;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
output 	Equal8;
input 	basic_reconfig_waitrequest2;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
input 	pll_go;
input 	uif_mode_0;
output 	Mux0;
output 	Mux3;
input 	WideOr0;
input 	pll_type;
input 	mif_rec_addr_7;
input 	mif_rec_addr_5;
input 	mif_rec_addr_6;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \inst_pll_ctrl|uif_rdata[3]~q ;
wire \inst_pll_ctrl|uif_rdata[4]~q ;
wire \inst_pll_ctrl|uif_rdata[5]~q ;
wire \inst_pll_ctrl|uif_rdata[6]~q ;
wire \inst_pll_ctrl|uif_rdata[7]~q ;
wire \inst_pll_ctrl|uif_rdata[8]~q ;
wire \inst_pll_ctrl|uif_rdata[9]~q ;
wire \inst_pll_ctrl|uif_rdata[10]~q ;
wire \inst_pll_ctrl|uif_rdata[11]~q ;
wire \inst_pll_ctrl|uif_rdata[12]~q ;
wire \inst_pll_ctrl|uif_rdata[13]~q ;
wire \inst_pll_ctrl|uif_rdata[14]~q ;
wire \inst_pll_ctrl|uif_rdata[15]~q ;
wire \inst_pll_ctrl|uif_rdata[16]~q ;
wire \inst_pll_ctrl|uif_rdata[17]~q ;
wire \inst_pll_ctrl|uif_rdata[18]~q ;
wire \inst_pll_ctrl|uif_rdata[19]~q ;
wire \inst_pll_ctrl|ctrl_wdata[1]~q ;
wire \inst_pll_ctrl|ctrl_addr[1]~q ;
wire \inst_pll_ctrl|ctrl_wdata[2]~q ;
wire \inst_pll_ctrl|ctrl_addr[5]~q ;
wire \inst_pll_ctrl|ctrl_wdata[0]~q ;
wire \inst_pll_ctrl|ctrl_addr[0]~q ;
wire \inst_pll_ctrl|ctrl_addr[4]~q ;
wire \inst_pll_ctrl|ctrl_wdata[5]~q ;
wire \inst_pll_ctrl|ctrl_wdata[9]~q ;
wire \inst_pll_ctrl|ctrl_wdata[13]~q ;
wire \inst_pll_ctrl|ctrl_wdata[14]~q ;
wire \inst_pll_ctrl|ctrl_wdata[15]~q ;
wire \inst_pll_uif|uif_writedata[0]~q ;
wire \inst_pll_uif|uif_mode[1]~q ;
wire \inst_pll_uif|uif_mode[0]~q ;
wire \inst_pll_ctrl|Equal4~0_combout ;
wire \inst_pll_ctrl|uif_rdata[0]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[0]~q ;
wire \inst_pll_uif|uif_addr_offset[0]~q ;
wire \inst_pll_uif|uif_writedata[1]~q ;
wire \inst_pll_ctrl|uif_rdata[1]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[1]~q ;
wire \inst_pll_uif|uif_addr_offset[1]~q ;
wire \inst_pll_uif|uif_writedata[2]~q ;
wire \inst_pll_ctrl|uif_rdata[2]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[2]~q ;
wire \inst_pll_uif|uif_addr_offset[2]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[3]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[4]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[5]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[6]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[7]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[8]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ;
wire \inst_pll_uif|uif_logical_ch_addr[9]~q ;
wire \inst_pll_ctrl|uif_addr_err~q ;
wire \inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ;
wire \inst_pll_ctrl|uif_rdata[20]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ;
wire \inst_pll_ctrl|uif_rdata[21]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ;
wire \inst_pll_ctrl|uif_rdata[22]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ;
wire \inst_pll_ctrl|uif_rdata[23]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ;
wire \inst_pll_ctrl|uif_rdata[24]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ;
wire \inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ;
wire \inst_pll_ctrl|ctrl_go~q ;
wire \inst_pll_ctrl|ctrl_lock~q ;
wire \inst_pll_ctrl|ctrl_opcode[2]~q ;
wire \inst_pll_ctrl|ctrl_opcode[0]~q ;
wire \inst_pll_uif|uif_go~q ;
wire \inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ;
wire \inst_pll_ctrl|ctrl_lch[4]~0_combout ;
wire \inst_pll_ctrl|ctrl_lch[5]~1_combout ;
wire \inst_pll_ctrl|ctrl_lch[2]~2_combout ;
wire \inst_pll_ctrl|ctrl_lch[3]~3_combout ;
wire \inst_pll_ctrl|ctrl_lch[0]~4_combout ;
wire \inst_pll_ctrl|ctrl_lch[1]~5_combout ;
wire \inst_pll_ctrl|ctrl_lch[8]~6_combout ;
wire \inst_pll_ctrl|ctrl_lch[9]~7_combout ;
wire \inst_pll_ctrl|ctrl_lch[6]~8_combout ;
wire \inst_pll_ctrl|ctrl_lch[7]~9_combout ;
wire \inst_pll_ctrl|ctrl_wdata[3]~q ;
wire \inst_pll_ctrl|ctrl_wdata[4]~q ;
wire \inst_pll_ctrl|ctrl_wdata[6]~q ;
wire \inst_pll_ctrl|ctrl_wdata[7]~q ;
wire \inst_pll_ctrl|ctrl_wdata[8]~q ;
wire \inst_pll_ctrl|ctrl_wdata[10]~q ;
wire \inst_pll_ctrl|ctrl_wdata[11]~q ;
wire \inst_pll_ctrl|ctrl_wdata[12]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ;
wire \inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ;


RECONFIGURE_IP_alt_xreconf_cif_2 inst_xreconf_cif(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.ctrl_wdata_1(\inst_pll_ctrl|ctrl_wdata[1]~q ),
	.ctrl_addr_1(\inst_pll_ctrl|ctrl_addr[1]~q ),
	.ctrl_wdata_2(\inst_pll_ctrl|ctrl_wdata[2]~q ),
	.ctrl_addr_5(\inst_pll_ctrl|ctrl_addr[5]~q ),
	.ctrl_wdata_0(\inst_pll_ctrl|ctrl_wdata[0]~q ),
	.ctrl_addr_0(\inst_pll_ctrl|ctrl_addr[0]~q ),
	.ctrl_addr_4(\inst_pll_ctrl|ctrl_addr[4]~q ),
	.ctrl_wdata_5(\inst_pll_ctrl|ctrl_wdata[5]~q ),
	.ctrl_wdata_9(\inst_pll_ctrl|ctrl_wdata[9]~q ),
	.ctrl_wdata_13(\inst_pll_ctrl|ctrl_wdata[13]~q ),
	.ctrl_wdata_14(\inst_pll_ctrl|ctrl_wdata[14]~q ),
	.ctrl_wdata_15(\inst_pll_ctrl|ctrl_wdata[15]~q ),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.master_write(master_write),
	.grant_8(grant_8),
	.mutex_req(mutex_req),
	.master_address_2(master_address_2),
	.master_address_0(master_address_0),
	.master_address_1(master_address_1),
	.lif_waitrequest(lif_waitrequest),
	.master_read(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.ph_readdata_0(\inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ),
	.ph_readdata_1(\inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ),
	.ph_readdata_2(\inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ),
	.ph_readdata_3(\inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ),
	.ph_readdata_4(\inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ),
	.ph_readdata_5(\inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ),
	.ph_readdata_6(\inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ),
	.ph_readdata_7(\inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ),
	.ph_readdata_8(\inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ),
	.ph_readdata_9(\inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ),
	.illegal_phy_ch(\inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ),
	.ph_readdata_10(\inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ),
	.ph_readdata_11(\inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ),
	.ph_readdata_12(\inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ),
	.ph_readdata_13(\inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ),
	.ph_readdata_14(\inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ),
	.ph_readdata_15(\inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ),
	.ph_readdata_16(\inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ),
	.ph_readdata_17(\inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ),
	.ph_readdata_18(\inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ),
	.ph_readdata_19(\inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ),
	.ph_readdata_20(\inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ),
	.ph_readdata_21(\inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ),
	.ph_readdata_22(\inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ),
	.ph_readdata_23(\inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ),
	.ph_readdata_24(\inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ),
	.ph_readdata_25(\inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ),
	.ph_readdata_26(\inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ),
	.ph_readdata_27(\inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ),
	.ph_readdata_28(\inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ),
	.ph_readdata_29(\inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ),
	.ph_readdata_30(\inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ),
	.ph_readdata_31(\inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ),
	.mutex_grant(mutex_grant),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.ctrl_go(\inst_pll_ctrl|ctrl_go~q ),
	.ctrl_lock(\inst_pll_ctrl|ctrl_lock~q ),
	.ctrl_opcode_2(\inst_pll_ctrl|ctrl_opcode[2]~q ),
	.ctrl_opcode_0(\inst_pll_ctrl|ctrl_opcode[0]~q ),
	.master_writedata_1(master_writedata_1),
	.master_writedata_2(master_writedata_2),
	.master_writedata_0(master_writedata_0),
	.master_writedata_3(master_writedata_3),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.master_writedata_11(master_writedata_11),
	.master_writedata_12(master_writedata_12),
	.master_writedata_13(master_writedata_13),
	.master_writedata_14(master_writedata_14),
	.master_writedata_15(master_writedata_15),
	.waitrequest_to_ctrl(\inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ),
	.ctrl_lch_4(\inst_pll_ctrl|ctrl_lch[4]~0_combout ),
	.ctrl_lch_5(\inst_pll_ctrl|ctrl_lch[5]~1_combout ),
	.ctrl_lch_2(\inst_pll_ctrl|ctrl_lch[2]~2_combout ),
	.ctrl_lch_3(\inst_pll_ctrl|ctrl_lch[3]~3_combout ),
	.ctrl_lch_0(\inst_pll_ctrl|ctrl_lch[0]~4_combout ),
	.ctrl_lch_1(\inst_pll_ctrl|ctrl_lch[1]~5_combout ),
	.ctrl_lch_8(\inst_pll_ctrl|ctrl_lch[8]~6_combout ),
	.ctrl_lch_9(\inst_pll_ctrl|ctrl_lch[9]~7_combout ),
	.ctrl_lch_6(\inst_pll_ctrl|ctrl_lch[6]~8_combout ),
	.ctrl_lch_7(\inst_pll_ctrl|ctrl_lch[7]~9_combout ),
	.ctrl_wdata_3(\inst_pll_ctrl|ctrl_wdata[3]~q ),
	.ctrl_wdata_4(\inst_pll_ctrl|ctrl_wdata[4]~q ),
	.ctrl_wdata_6(\inst_pll_ctrl|ctrl_wdata[6]~q ),
	.ctrl_wdata_7(\inst_pll_ctrl|ctrl_wdata[7]~q ),
	.ctrl_wdata_8(\inst_pll_ctrl|ctrl_wdata[8]~q ),
	.ctrl_wdata_10(\inst_pll_ctrl|ctrl_wdata[10]~q ),
	.ctrl_wdata_11(\inst_pll_ctrl|ctrl_wdata[11]~q ),
	.ctrl_wdata_12(\inst_pll_ctrl|ctrl_wdata[12]~q ),
	.readdata_for_user_0(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q ),
	.readdata_for_user_1(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ),
	.readdata_for_user_2(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ),
	.readdata_for_user_3(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ),
	.readdata_for_user_4(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ),
	.readdata_for_user_5(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ),
	.readdata_for_user_6(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ),
	.readdata_for_user_7(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ),
	.readdata_for_user_8(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ),
	.readdata_for_user_9(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ),
	.readdata_for_user_10(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ),
	.readdata_for_user_11(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ),
	.readdata_for_user_12(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ),
	.readdata_for_user_13(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ),
	.readdata_for_user_14(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ),
	.readdata_for_user_15(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ),
	.readdata_for_user_16(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ),
	.readdata_for_user_17(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ),
	.readdata_for_user_18(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ),
	.readdata_for_user_19(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ),
	.readdata_for_user_20(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.readdata_for_user_21(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.readdata_for_user_22(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.readdata_for_user_23(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.readdata_for_user_24(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.mgmt_clk_clk(mgmt_clk_clk));

RECONFIGURE_IP_av_xcvr_reconfig_pll_ctrl inst_pll_ctrl(
	.uif_rdata_3(\inst_pll_ctrl|uif_rdata[3]~q ),
	.uif_rdata_4(\inst_pll_ctrl|uif_rdata[4]~q ),
	.uif_rdata_5(\inst_pll_ctrl|uif_rdata[5]~q ),
	.uif_rdata_6(\inst_pll_ctrl|uif_rdata[6]~q ),
	.uif_rdata_7(\inst_pll_ctrl|uif_rdata[7]~q ),
	.uif_rdata_8(\inst_pll_ctrl|uif_rdata[8]~q ),
	.uif_rdata_9(\inst_pll_ctrl|uif_rdata[9]~q ),
	.uif_rdata_10(\inst_pll_ctrl|uif_rdata[10]~q ),
	.uif_rdata_11(\inst_pll_ctrl|uif_rdata[11]~q ),
	.uif_rdata_12(\inst_pll_ctrl|uif_rdata[12]~q ),
	.uif_rdata_13(\inst_pll_ctrl|uif_rdata[13]~q ),
	.uif_rdata_14(\inst_pll_ctrl|uif_rdata[14]~q ),
	.uif_rdata_15(\inst_pll_ctrl|uif_rdata[15]~q ),
	.uif_rdata_16(\inst_pll_ctrl|uif_rdata[16]~q ),
	.uif_rdata_17(\inst_pll_ctrl|uif_rdata[17]~q ),
	.uif_rdata_18(\inst_pll_ctrl|uif_rdata[18]~q ),
	.uif_rdata_19(\inst_pll_ctrl|uif_rdata[19]~q ),
	.ctrl_wdata_1(\inst_pll_ctrl|ctrl_wdata[1]~q ),
	.ctrl_addr_1(\inst_pll_ctrl|ctrl_addr[1]~q ),
	.ctrl_wdata_2(\inst_pll_ctrl|ctrl_wdata[2]~q ),
	.ctrl_addr_5(\inst_pll_ctrl|ctrl_addr[5]~q ),
	.ctrl_wdata_0(\inst_pll_ctrl|ctrl_wdata[0]~q ),
	.ctrl_addr_0(\inst_pll_ctrl|ctrl_addr[0]~q ),
	.ctrl_addr_4(\inst_pll_ctrl|ctrl_addr[4]~q ),
	.ctrl_wdata_5(\inst_pll_ctrl|ctrl_wdata[5]~q ),
	.ctrl_wdata_9(\inst_pll_ctrl|ctrl_wdata[9]~q ),
	.ctrl_wdata_13(\inst_pll_ctrl|ctrl_wdata[13]~q ),
	.ctrl_wdata_14(\inst_pll_ctrl|ctrl_wdata[14]~q ),
	.ctrl_wdata_15(\inst_pll_ctrl|ctrl_wdata[15]~q ),
	.pll_mif_busy1(pll_mif_busy),
	.reset(ifsel_notdone_resync),
	.uif_logical_ch_addr_0(uif_logical_ch_addr_0),
	.uif_wdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\inst_pll_uif|uif_writedata[2]~q ,\inst_pll_uif|uif_writedata[1]~q ,\inst_pll_uif|uif_writedata[0]~q }),
	.uif_mode_1(\inst_pll_uif|uif_mode[1]~q ),
	.uif_mode_0(\inst_pll_uif|uif_mode[0]~q ),
	.Equal4(\inst_pll_ctrl|Equal4~0_combout ),
	.uif_rdata_0(\inst_pll_ctrl|uif_rdata[0]~q ),
	.uif_logical_ch_addr_01(\inst_pll_uif|uif_logical_ch_addr[0]~q ),
	.uif_addr_offset_0(\inst_pll_uif|uif_addr_offset[0]~q ),
	.uif_logical_ch_addr_1(uif_logical_ch_addr_1),
	.uif_rdata_1(\inst_pll_ctrl|uif_rdata[1]~q ),
	.uif_logical_ch_addr_11(\inst_pll_uif|uif_logical_ch_addr[1]~q ),
	.uif_addr_offset_1(\inst_pll_uif|uif_addr_offset[1]~q ),
	.uif_logical_ch_addr_2(uif_logical_ch_addr_2),
	.uif_rdata_2(\inst_pll_ctrl|uif_rdata[2]~q ),
	.uif_logical_ch_addr_21(\inst_pll_uif|uif_logical_ch_addr[2]~q ),
	.uif_addr_offset_2(\inst_pll_uif|uif_addr_offset[2]~q ),
	.uif_logical_ch_addr_3(uif_logical_ch_addr_3),
	.uif_logical_ch_addr_31(\inst_pll_uif|uif_logical_ch_addr[3]~q ),
	.uif_logical_ch_addr_4(uif_logical_ch_addr_4),
	.uif_logical_ch_addr_41(\inst_pll_uif|uif_logical_ch_addr[4]~q ),
	.uif_logical_ch_addr_5(uif_logical_ch_addr_5),
	.uif_logical_ch_addr_51(\inst_pll_uif|uif_logical_ch_addr[5]~q ),
	.uif_logical_ch_addr_6(uif_logical_ch_addr_6),
	.uif_logical_ch_addr_61(\inst_pll_uif|uif_logical_ch_addr[6]~q ),
	.uif_logical_ch_addr_7(uif_logical_ch_addr_7),
	.uif_logical_ch_addr_71(\inst_pll_uif|uif_logical_ch_addr[7]~q ),
	.uif_logical_ch_addr_8(\inst_pll_uif|uif_logical_ch_addr[8]~q ),
	.uif_logical_ch_addr_81(uif_logical_ch_addr_8),
	.uif_logical_ch_addr_9(uif_logical_ch_addr_9),
	.uif_logical_ch_addr_91(\inst_pll_uif|uif_logical_ch_addr[9]~q ),
	.uif_addr_err1(\inst_pll_ctrl|uif_addr_err~q ),
	.uif_rdata_20(\inst_pll_ctrl|uif_rdata[20]~q ),
	.uif_rdata_21(\inst_pll_ctrl|uif_rdata[21]~q ),
	.uif_rdata_22(\inst_pll_ctrl|uif_rdata[22]~q ),
	.uif_rdata_23(\inst_pll_ctrl|uif_rdata[23]~q ),
	.uif_rdata_24(\inst_pll_ctrl|uif_rdata[24]~q ),
	.ctrl_go1(\inst_pll_ctrl|ctrl_go~q ),
	.ctrl_lock1(\inst_pll_ctrl|ctrl_lock~q ),
	.ctrl_opcode_2(\inst_pll_ctrl|ctrl_opcode[2]~q ),
	.ctrl_opcode_0(\inst_pll_ctrl|ctrl_opcode[0]~q ),
	.pll_go(pll_go),
	.uif_go(\inst_pll_uif|uif_go~q ),
	.waitrequest_to_ctrl(\inst_xreconf_cif|inst_basic_acq|waitrequest_to_ctrl~q ),
	.ctrl_lch_4(\inst_pll_ctrl|ctrl_lch[4]~0_combout ),
	.ctrl_lch_5(\inst_pll_ctrl|ctrl_lch[5]~1_combout ),
	.ctrl_lch_2(\inst_pll_ctrl|ctrl_lch[2]~2_combout ),
	.ctrl_lch_3(\inst_pll_ctrl|ctrl_lch[3]~3_combout ),
	.ctrl_lch_0(\inst_pll_ctrl|ctrl_lch[0]~4_combout ),
	.ctrl_lch_1(\inst_pll_ctrl|ctrl_lch[1]~5_combout ),
	.ctrl_lch_8(\inst_pll_ctrl|ctrl_lch[8]~6_combout ),
	.ctrl_lch_9(\inst_pll_ctrl|ctrl_lch[9]~7_combout ),
	.ctrl_lch_6(\inst_pll_ctrl|ctrl_lch[6]~8_combout ),
	.ctrl_lch_7(\inst_pll_ctrl|ctrl_lch[7]~9_combout ),
	.ctrl_wdata_3(\inst_pll_ctrl|ctrl_wdata[3]~q ),
	.ctrl_wdata_4(\inst_pll_ctrl|ctrl_wdata[4]~q ),
	.ctrl_wdata_6(\inst_pll_ctrl|ctrl_wdata[6]~q ),
	.ctrl_wdata_7(\inst_pll_ctrl|ctrl_wdata[7]~q ),
	.ctrl_wdata_8(\inst_pll_ctrl|ctrl_wdata[8]~q ),
	.ctrl_wdata_10(\inst_pll_ctrl|ctrl_wdata[10]~q ),
	.ctrl_wdata_11(\inst_pll_ctrl|ctrl_wdata[11]~q ),
	.ctrl_wdata_12(\inst_pll_ctrl|ctrl_wdata[12]~q ),
	.ctrl_rdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[19]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[18]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[17]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[16]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[15]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[14]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[13]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[12]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[11]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[10]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[9]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[8]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[7]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[6]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[5]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[4]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[3]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[2]~q ,\inst_xreconf_cif|inst_basic_acq|readdata_for_user[1]~q ,
\inst_xreconf_cif|inst_basic_acq|readdata_for_user[0]~q }),
	.pll_type(pll_type),
	.readdata_for_user_20(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[20]~q ),
	.readdata_for_user_21(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[21]~q ),
	.readdata_for_user_22(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[22]~q ),
	.readdata_for_user_23(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[23]~q ),
	.readdata_for_user_24(\inst_xreconf_cif|inst_basic_acq|readdata_for_user[24]~q ),
	.mif_rec_addr_7(mif_rec_addr_7),
	.mif_rec_addr_5(mif_rec_addr_5),
	.mif_rec_addr_6(mif_rec_addr_6),
	.clk(mgmt_clk_clk));

RECONFIGURE_IP_alt_xreconf_uif_2 inst_pll_uif(
	.user_reconfig_readdata_10(user_reconfig_readdata_10),
	.user_reconfig_readdata_11(user_reconfig_readdata_11),
	.user_reconfig_readdata_12(user_reconfig_readdata_12),
	.user_reconfig_readdata_13(user_reconfig_readdata_13),
	.user_reconfig_readdata_14(user_reconfig_readdata_14),
	.user_reconfig_readdata_15(user_reconfig_readdata_15),
	.user_reconfig_readdata_16(user_reconfig_readdata_16),
	.user_reconfig_readdata_17(user_reconfig_readdata_17),
	.user_reconfig_readdata_18(user_reconfig_readdata_18),
	.user_reconfig_readdata_19(user_reconfig_readdata_19),
	.user_reconfig_readdata_20(user_reconfig_readdata_20),
	.user_reconfig_readdata_21(user_reconfig_readdata_21),
	.user_reconfig_readdata_22(user_reconfig_readdata_22),
	.user_reconfig_readdata_23(user_reconfig_readdata_23),
	.user_reconfig_readdata_24(user_reconfig_readdata_24),
	.uif_rdata_3(\inst_pll_ctrl|uif_rdata[3]~q ),
	.uif_rdata_4(\inst_pll_ctrl|uif_rdata[4]~q ),
	.uif_rdata_5(\inst_pll_ctrl|uif_rdata[5]~q ),
	.uif_rdata_6(\inst_pll_ctrl|uif_rdata[6]~q ),
	.uif_rdata_7(\inst_pll_ctrl|uif_rdata[7]~q ),
	.uif_rdata_8(\inst_pll_ctrl|uif_rdata[8]~q ),
	.uif_rdata_9(\inst_pll_ctrl|uif_rdata[9]~q ),
	.uif_rdata_10(\inst_pll_ctrl|uif_rdata[10]~q ),
	.uif_rdata_11(\inst_pll_ctrl|uif_rdata[11]~q ),
	.uif_rdata_12(\inst_pll_ctrl|uif_rdata[12]~q ),
	.uif_rdata_13(\inst_pll_ctrl|uif_rdata[13]~q ),
	.uif_rdata_14(\inst_pll_ctrl|uif_rdata[14]~q ),
	.uif_rdata_15(\inst_pll_ctrl|uif_rdata[15]~q ),
	.uif_rdata_16(\inst_pll_ctrl|uif_rdata[16]~q ),
	.uif_rdata_17(\inst_pll_ctrl|uif_rdata[17]~q ),
	.uif_rdata_18(\inst_pll_ctrl|uif_rdata[18]~q ),
	.uif_rdata_19(\inst_pll_ctrl|uif_rdata[19]~q ),
	.user_reconfig_readdata_0(user_reconfig_readdata_0),
	.Equal4(Equal4),
	.user_reconfig_readdata_1(user_reconfig_readdata_1),
	.user_reconfig_readdata_2(user_reconfig_readdata_2),
	.user_reconfig_readdata_3(user_reconfig_readdata_3),
	.user_reconfig_readdata_4(user_reconfig_readdata_4),
	.user_reconfig_readdata_5(user_reconfig_readdata_5),
	.user_reconfig_readdata_6(user_reconfig_readdata_6),
	.user_reconfig_readdata_7(user_reconfig_readdata_7),
	.user_reconfig_readdata_8(user_reconfig_readdata_8),
	.user_reconfig_readdata_9(user_reconfig_readdata_9),
	.user_reconfig_readdata_25(user_reconfig_readdata_25),
	.user_reconfig_readdata_26(user_reconfig_readdata_26),
	.user_reconfig_readdata_27(user_reconfig_readdata_27),
	.user_reconfig_readdata_28(user_reconfig_readdata_28),
	.user_reconfig_readdata_29(user_reconfig_readdata_29),
	.user_reconfig_readdata_30(user_reconfig_readdata_30),
	.user_reconfig_readdata_31(user_reconfig_readdata_31),
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg(launch_reg),
	.wait_reg(wait_reg),
	.pll_mif_busy(pll_mif_busy),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.uif_writedata_0(\inst_pll_uif|uif_writedata[0]~q ),
	.uif_mode_1(\inst_pll_uif|uif_mode[1]~q ),
	.uif_mode_0(\inst_pll_uif|uif_mode[0]~q ),
	.Equal41(\inst_pll_ctrl|Equal4~0_combout ),
	.uif_rdata_0(\inst_pll_ctrl|uif_rdata[0]~q ),
	.ph_readdata_0(\inst_xreconf_cif|inst_basic_acq|ph_readdata[0]~q ),
	.uif_logical_ch_addr_0(\inst_pll_uif|uif_logical_ch_addr[0]~q ),
	.uif_addr_offset_0(\inst_pll_uif|uif_addr_offset[0]~q ),
	.comb(comb),
	.uif_writedata_1(\inst_pll_uif|uif_writedata[1]~q ),
	.uif_rdata_1(\inst_pll_ctrl|uif_rdata[1]~q ),
	.ph_readdata_1(\inst_xreconf_cif|inst_basic_acq|ph_readdata[1]~q ),
	.uif_logical_ch_addr_1(\inst_pll_uif|uif_logical_ch_addr[1]~q ),
	.uif_addr_offset_1(\inst_pll_uif|uif_addr_offset[1]~q ),
	.uif_writedata_2(\inst_pll_uif|uif_writedata[2]~q ),
	.uif_rdata_2(\inst_pll_ctrl|uif_rdata[2]~q ),
	.ph_readdata_2(\inst_xreconf_cif|inst_basic_acq|ph_readdata[2]~q ),
	.uif_logical_ch_addr_2(\inst_pll_uif|uif_logical_ch_addr[2]~q ),
	.uif_addr_offset_2(\inst_pll_uif|uif_addr_offset[2]~q ),
	.ph_readdata_3(\inst_xreconf_cif|inst_basic_acq|ph_readdata[3]~q ),
	.uif_logical_ch_addr_3(\inst_pll_uif|uif_logical_ch_addr[3]~q ),
	.user_reconfig_readdata_101(user_reconfig_readdata_101),
	.ph_readdata_4(\inst_xreconf_cif|inst_basic_acq|ph_readdata[4]~q ),
	.uif_logical_ch_addr_4(\inst_pll_uif|uif_logical_ch_addr[4]~q ),
	.ph_readdata_5(\inst_xreconf_cif|inst_basic_acq|ph_readdata[5]~q ),
	.uif_logical_ch_addr_5(\inst_pll_uif|uif_logical_ch_addr[5]~q ),
	.ph_readdata_6(\inst_xreconf_cif|inst_basic_acq|ph_readdata[6]~q ),
	.uif_logical_ch_addr_6(\inst_pll_uif|uif_logical_ch_addr[6]~q ),
	.ph_readdata_7(\inst_xreconf_cif|inst_basic_acq|ph_readdata[7]~q ),
	.uif_logical_ch_addr_7(\inst_pll_uif|uif_logical_ch_addr[7]~q ),
	.uif_logical_ch_addr_8(\inst_pll_uif|uif_logical_ch_addr[8]~q ),
	.ph_readdata_8(\inst_xreconf_cif|inst_basic_acq|ph_readdata[8]~q ),
	.ph_readdata_9(\inst_xreconf_cif|inst_basic_acq|ph_readdata[9]~q ),
	.uif_logical_ch_addr_9(\inst_pll_uif|uif_logical_ch_addr[9]~q ),
	.uif_addr_err(\inst_pll_ctrl|uif_addr_err~q ),
	.illegal_phy_ch(\inst_xreconf_cif|inst_basic_acq|illegal_phy_ch~q ),
	.ph_readdata_10(\inst_xreconf_cif|inst_basic_acq|ph_readdata[10]~q ),
	.ph_readdata_11(\inst_xreconf_cif|inst_basic_acq|ph_readdata[11]~q ),
	.ph_readdata_12(\inst_xreconf_cif|inst_basic_acq|ph_readdata[12]~q ),
	.ph_readdata_13(\inst_xreconf_cif|inst_basic_acq|ph_readdata[13]~q ),
	.ph_readdata_14(\inst_xreconf_cif|inst_basic_acq|ph_readdata[14]~q ),
	.ph_readdata_15(\inst_xreconf_cif|inst_basic_acq|ph_readdata[15]~q ),
	.ph_readdata_16(\inst_xreconf_cif|inst_basic_acq|ph_readdata[16]~q ),
	.ph_readdata_17(\inst_xreconf_cif|inst_basic_acq|ph_readdata[17]~q ),
	.ph_readdata_18(\inst_xreconf_cif|inst_basic_acq|ph_readdata[18]~q ),
	.ph_readdata_19(\inst_xreconf_cif|inst_basic_acq|ph_readdata[19]~q ),
	.ph_readdata_20(\inst_xreconf_cif|inst_basic_acq|ph_readdata[20]~q ),
	.uif_rdata_20(\inst_pll_ctrl|uif_rdata[20]~q ),
	.ph_readdata_21(\inst_xreconf_cif|inst_basic_acq|ph_readdata[21]~q ),
	.uif_rdata_21(\inst_pll_ctrl|uif_rdata[21]~q ),
	.ph_readdata_22(\inst_xreconf_cif|inst_basic_acq|ph_readdata[22]~q ),
	.uif_rdata_22(\inst_pll_ctrl|uif_rdata[22]~q ),
	.ph_readdata_23(\inst_xreconf_cif|inst_basic_acq|ph_readdata[23]~q ),
	.uif_rdata_23(\inst_pll_ctrl|uif_rdata[23]~q ),
	.ph_readdata_24(\inst_xreconf_cif|inst_basic_acq|ph_readdata[24]~q ),
	.uif_rdata_24(\inst_pll_ctrl|uif_rdata[24]~q ),
	.ph_readdata_25(\inst_xreconf_cif|inst_basic_acq|ph_readdata[25]~q ),
	.ph_readdata_26(\inst_xreconf_cif|inst_basic_acq|ph_readdata[26]~q ),
	.ph_readdata_27(\inst_xreconf_cif|inst_basic_acq|ph_readdata[27]~q ),
	.ph_readdata_28(\inst_xreconf_cif|inst_basic_acq|ph_readdata[28]~q ),
	.ph_readdata_29(\inst_xreconf_cif|inst_basic_acq|ph_readdata[29]~q ),
	.ph_readdata_30(\inst_xreconf_cif|inst_basic_acq|ph_readdata[30]~q ),
	.ph_readdata_31(\inst_xreconf_cif|inst_basic_acq|ph_readdata[31]~q ),
	.uif_go1(\inst_pll_uif|uif_go~q ),
	.uif_mode_01(uif_mode_0),
	.Mux0(Mux0),
	.Mux3(Mux3),
	.WideOr0(WideOr0),
	.reconfig_mgmt_address_1(reconfig_mgmt_address_1),
	.reconfig_mgmt_address_0(reconfig_mgmt_address_0),
	.reconfig_mgmt_address_2(reconfig_mgmt_address_2),
	.reconfig_mgmt_write(reconfig_mgmt_write),
	.reconfig_mgmt_read(reconfig_mgmt_read),
	.mgmt_clk_clk(mgmt_clk_clk),
	.reconfig_mgmt_writedata_0(reconfig_mgmt_writedata_0),
	.reconfig_mgmt_writedata_1(reconfig_mgmt_writedata_1),
	.reconfig_mgmt_writedata_2(reconfig_mgmt_writedata_2),
	.reconfig_mgmt_writedata_3(reconfig_mgmt_writedata_3),
	.reconfig_mgmt_writedata_16(reconfig_mgmt_writedata_16),
	.reconfig_mgmt_writedata_17(reconfig_mgmt_writedata_17),
	.reconfig_mgmt_writedata_18(reconfig_mgmt_writedata_18),
	.reconfig_mgmt_writedata_19(reconfig_mgmt_writedata_19),
	.reconfig_mgmt_writedata_20(reconfig_mgmt_writedata_20),
	.reconfig_mgmt_writedata_4(reconfig_mgmt_writedata_4),
	.reconfig_mgmt_writedata_21(reconfig_mgmt_writedata_21),
	.reconfig_mgmt_writedata_5(reconfig_mgmt_writedata_5),
	.reconfig_mgmt_writedata_22(reconfig_mgmt_writedata_22),
	.reconfig_mgmt_writedata_6(reconfig_mgmt_writedata_6),
	.reconfig_mgmt_writedata_23(reconfig_mgmt_writedata_23),
	.reconfig_mgmt_writedata_7(reconfig_mgmt_writedata_7),
	.reconfig_mgmt_writedata_24(reconfig_mgmt_writedata_24),
	.reconfig_mgmt_writedata_8(reconfig_mgmt_writedata_8),
	.reconfig_mgmt_writedata_25(reconfig_mgmt_writedata_25),
	.reconfig_mgmt_writedata_9(reconfig_mgmt_writedata_9),
	.reconfig_mgmt_writedata_26(reconfig_mgmt_writedata_26),
	.reconfig_mgmt_writedata_10(reconfig_mgmt_writedata_10),
	.reconfig_mgmt_writedata_27(reconfig_mgmt_writedata_27),
	.reconfig_mgmt_writedata_11(reconfig_mgmt_writedata_11),
	.reconfig_mgmt_writedata_28(reconfig_mgmt_writedata_28),
	.reconfig_mgmt_writedata_12(reconfig_mgmt_writedata_12),
	.reconfig_mgmt_writedata_29(reconfig_mgmt_writedata_29),
	.reconfig_mgmt_writedata_13(reconfig_mgmt_writedata_13),
	.reconfig_mgmt_writedata_30(reconfig_mgmt_writedata_30),
	.reconfig_mgmt_writedata_14(reconfig_mgmt_writedata_14),
	.reconfig_mgmt_writedata_31(reconfig_mgmt_writedata_31),
	.reconfig_mgmt_writedata_15(reconfig_mgmt_writedata_15));

endmodule

module RECONFIGURE_IP_alt_xreconf_cif_2 (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	ctrl_wdata_1,
	ctrl_addr_1,
	ctrl_wdata_2,
	ctrl_addr_5,
	ctrl_wdata_0,
	ctrl_addr_0,
	ctrl_addr_4,
	ctrl_wdata_5,
	ctrl_wdata_9,
	ctrl_wdata_13,
	ctrl_wdata_14,
	ctrl_wdata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write,
	grant_8,
	mutex_req,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	ifsel_notdone_resync,
	ph_readdata_0,
	ph_readdata_1,
	ph_readdata_2,
	ph_readdata_3,
	ph_readdata_4,
	ph_readdata_5,
	ph_readdata_6,
	ph_readdata_7,
	ph_readdata_8,
	ph_readdata_9,
	illegal_phy_ch,
	ph_readdata_10,
	ph_readdata_11,
	ph_readdata_12,
	ph_readdata_13,
	ph_readdata_14,
	ph_readdata_15,
	ph_readdata_16,
	ph_readdata_17,
	ph_readdata_18,
	ph_readdata_19,
	ph_readdata_20,
	ph_readdata_21,
	ph_readdata_22,
	ph_readdata_23,
	ph_readdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	mutex_grant,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	ctrl_go,
	ctrl_lock,
	ctrl_opcode_2,
	ctrl_opcode_0,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	waitrequest_to_ctrl,
	ctrl_lch_4,
	ctrl_lch_5,
	ctrl_lch_2,
	ctrl_lch_3,
	ctrl_lch_0,
	ctrl_lch_1,
	ctrl_lch_8,
	ctrl_lch_9,
	ctrl_lch_6,
	ctrl_lch_7,
	ctrl_wdata_3,
	ctrl_wdata_4,
	ctrl_wdata_6,
	ctrl_wdata_7,
	ctrl_wdata_8,
	ctrl_wdata_10,
	ctrl_wdata_11,
	ctrl_wdata_12,
	readdata_for_user_0,
	readdata_for_user_1,
	readdata_for_user_2,
	readdata_for_user_3,
	readdata_for_user_4,
	readdata_for_user_5,
	readdata_for_user_6,
	readdata_for_user_7,
	readdata_for_user_8,
	readdata_for_user_9,
	readdata_for_user_10,
	readdata_for_user_11,
	readdata_for_user_12,
	readdata_for_user_13,
	readdata_for_user_14,
	readdata_for_user_15,
	readdata_for_user_16,
	readdata_for_user_17,
	readdata_for_user_18,
	readdata_for_user_19,
	readdata_for_user_20,
	readdata_for_user_21,
	readdata_for_user_22,
	readdata_for_user_23,
	readdata_for_user_24,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_16;
input 	basic_reconfig_readdata_17;
input 	basic_reconfig_readdata_18;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
input 	ctrl_wdata_1;
input 	ctrl_addr_1;
input 	ctrl_wdata_2;
input 	ctrl_addr_5;
input 	ctrl_wdata_0;
input 	ctrl_addr_0;
input 	ctrl_addr_4;
input 	ctrl_wdata_5;
input 	ctrl_wdata_9;
input 	ctrl_wdata_13;
input 	ctrl_wdata_14;
input 	ctrl_wdata_15;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write;
input 	grant_8;
output 	mutex_req;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	ifsel_notdone_resync;
output 	ph_readdata_0;
output 	ph_readdata_1;
output 	ph_readdata_2;
output 	ph_readdata_3;
output 	ph_readdata_4;
output 	ph_readdata_5;
output 	ph_readdata_6;
output 	ph_readdata_7;
output 	ph_readdata_8;
output 	ph_readdata_9;
output 	illegal_phy_ch;
output 	ph_readdata_10;
output 	ph_readdata_11;
output 	ph_readdata_12;
output 	ph_readdata_13;
output 	ph_readdata_14;
output 	ph_readdata_15;
output 	ph_readdata_16;
output 	ph_readdata_17;
output 	ph_readdata_18;
output 	ph_readdata_19;
output 	ph_readdata_20;
output 	ph_readdata_21;
output 	ph_readdata_22;
output 	ph_readdata_23;
output 	ph_readdata_24;
output 	ph_readdata_25;
output 	ph_readdata_26;
output 	ph_readdata_27;
output 	ph_readdata_28;
output 	ph_readdata_29;
output 	ph_readdata_30;
output 	ph_readdata_31;
output 	mutex_grant;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
output 	Equal8;
input 	basic_reconfig_waitrequest2;
input 	ctrl_go;
input 	ctrl_lock;
input 	ctrl_opcode_2;
input 	ctrl_opcode_0;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
output 	waitrequest_to_ctrl;
input 	ctrl_lch_4;
input 	ctrl_lch_5;
input 	ctrl_lch_2;
input 	ctrl_lch_3;
input 	ctrl_lch_0;
input 	ctrl_lch_1;
input 	ctrl_lch_8;
input 	ctrl_lch_9;
input 	ctrl_lch_6;
input 	ctrl_lch_7;
input 	ctrl_wdata_3;
input 	ctrl_wdata_4;
input 	ctrl_wdata_6;
input 	ctrl_wdata_7;
input 	ctrl_wdata_8;
input 	ctrl_wdata_10;
input 	ctrl_wdata_11;
input 	ctrl_wdata_12;
output 	readdata_for_user_0;
output 	readdata_for_user_1;
output 	readdata_for_user_2;
output 	readdata_for_user_3;
output 	readdata_for_user_4;
output 	readdata_for_user_5;
output 	readdata_for_user_6;
output 	readdata_for_user_7;
output 	readdata_for_user_8;
output 	readdata_for_user_9;
output 	readdata_for_user_10;
output 	readdata_for_user_11;
output 	readdata_for_user_12;
output 	readdata_for_user_13;
output 	readdata_for_user_14;
output 	readdata_for_user_15;
output 	readdata_for_user_16;
output 	readdata_for_user_17;
output 	readdata_for_user_18;
output 	readdata_for_user_19;
output 	readdata_for_user_20;
output 	readdata_for_user_21;
output 	readdata_for_user_22;
output 	readdata_for_user_23;
output 	readdata_for_user_24;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \inst_basic_acq|master_address[2]~q ;
wire \inst_basic_acq|master_address[1]~q ;
wire \inst_basic_acq|master_writedata[1]~q ;
wire \inst_basic_acq|master_writedata[2]~q ;
wire \inst_basic_acq|master_writedata[0]~q ;
wire \inst_basic_acq|master_writedata[3]~q ;


RECONFIGURE_IP_alt_arbiter_acq_4 mutex_inst(
	.grant_8(grant_8),
	.mutex_req(mutex_req),
	.master_address_2(\inst_basic_acq|master_address[2]~q ),
	.master_address_21(master_address_2),
	.master_address_1(\inst_basic_acq|master_address[1]~q ),
	.master_address_11(master_address_1),
	.mutex_grant1(mutex_grant),
	.master_writedata_1(\inst_basic_acq|master_writedata[1]~q ),
	.master_writedata_11(master_writedata_1),
	.master_writedata_2(\inst_basic_acq|master_writedata[2]~q ),
	.master_writedata_21(master_writedata_2),
	.master_writedata_0(\inst_basic_acq|master_writedata[0]~q ),
	.master_writedata_01(master_writedata_0),
	.master_writedata_3(\inst_basic_acq|master_writedata[3]~q ),
	.master_writedata_31(master_writedata_3));

RECONFIGURE_IP_alt_xreconf_basic_acq_2 inst_basic_acq(
	.basic_reconfig_readdata_12(basic_reconfig_readdata_12),
	.basic_reconfig_readdata_13(basic_reconfig_readdata_13),
	.basic_reconfig_readdata_14(basic_reconfig_readdata_14),
	.basic_reconfig_readdata_15(basic_reconfig_readdata_15),
	.basic_reconfig_readdata_16(basic_reconfig_readdata_16),
	.basic_reconfig_readdata_17(basic_reconfig_readdata_17),
	.basic_reconfig_readdata_18(basic_reconfig_readdata_18),
	.basic_reconfig_readdata_19(basic_reconfig_readdata_19),
	.basic_reconfig_readdata_20(basic_reconfig_readdata_20),
	.basic_reconfig_readdata_21(basic_reconfig_readdata_21),
	.basic_reconfig_readdata_22(basic_reconfig_readdata_22),
	.basic_reconfig_readdata_23(basic_reconfig_readdata_23),
	.basic_reconfig_readdata_24(basic_reconfig_readdata_24),
	.basic_reconfig_readdata_25(basic_reconfig_readdata_25),
	.basic_reconfig_readdata_26(basic_reconfig_readdata_26),
	.basic_reconfig_readdata_27(basic_reconfig_readdata_27),
	.basic_reconfig_readdata_28(basic_reconfig_readdata_28),
	.basic_reconfig_readdata_29(basic_reconfig_readdata_29),
	.basic_reconfig_readdata_30(basic_reconfig_readdata_30),
	.basic_reconfig_readdata_31(basic_reconfig_readdata_31),
	.ctrl_wdata_1(ctrl_wdata_1),
	.ctrl_addr_1(ctrl_addr_1),
	.ctrl_wdata_2(ctrl_wdata_2),
	.ctrl_addr_5(ctrl_addr_5),
	.ctrl_wdata_0(ctrl_wdata_0),
	.ctrl_addr_0(ctrl_addr_0),
	.ctrl_addr_4(ctrl_addr_4),
	.ctrl_wdata_5(ctrl_wdata_5),
	.ctrl_wdata_9(ctrl_wdata_9),
	.ctrl_wdata_13(ctrl_wdata_13),
	.ctrl_wdata_14(ctrl_wdata_14),
	.ctrl_wdata_15(ctrl_wdata_15),
	.basic_reconfig_readdata_0(basic_reconfig_readdata_0),
	.basic_reconfig_readdata_1(basic_reconfig_readdata_1),
	.basic_reconfig_readdata_2(basic_reconfig_readdata_2),
	.basic_reconfig_readdata_3(basic_reconfig_readdata_3),
	.basic_reconfig_readdata_4(basic_reconfig_readdata_4),
	.basic_reconfig_readdata_5(basic_reconfig_readdata_5),
	.basic_reconfig_readdata_6(basic_reconfig_readdata_6),
	.basic_reconfig_readdata_7(basic_reconfig_readdata_7),
	.basic_reconfig_readdata_8(basic_reconfig_readdata_8),
	.basic_reconfig_readdata_9(basic_reconfig_readdata_9),
	.basic_reconfig_readdata_10(basic_reconfig_readdata_10),
	.basic_reconfig_readdata_11(basic_reconfig_readdata_11),
	.master_write1(master_write),
	.mutex_req1(mutex_req),
	.master_address_2(\inst_basic_acq|master_address[2]~q ),
	.master_address_0(master_address_0),
	.master_address_1(\inst_basic_acq|master_address[1]~q ),
	.lif_waitrequest(lif_waitrequest),
	.master_read1(master_read),
	.basic_reconfig_waitrequest(basic_reconfig_waitrequest),
	.basic_reconfig_waitrequest1(basic_reconfig_waitrequest1),
	.reset(ifsel_notdone_resync),
	.ph_readdata_0(ph_readdata_0),
	.ph_readdata_1(ph_readdata_1),
	.ph_readdata_2(ph_readdata_2),
	.ph_readdata_3(ph_readdata_3),
	.ph_readdata_4(ph_readdata_4),
	.ph_readdata_5(ph_readdata_5),
	.ph_readdata_6(ph_readdata_6),
	.ph_readdata_7(ph_readdata_7),
	.ph_readdata_8(ph_readdata_8),
	.ph_readdata_9(ph_readdata_9),
	.illegal_phy_ch1(illegal_phy_ch),
	.ph_readdata_10(ph_readdata_10),
	.ph_readdata_11(ph_readdata_11),
	.ph_readdata_12(ph_readdata_12),
	.ph_readdata_13(ph_readdata_13),
	.ph_readdata_14(ph_readdata_14),
	.ph_readdata_15(ph_readdata_15),
	.ph_readdata_16(ph_readdata_16),
	.ph_readdata_17(ph_readdata_17),
	.ph_readdata_18(ph_readdata_18),
	.ph_readdata_19(ph_readdata_19),
	.ph_readdata_20(ph_readdata_20),
	.ph_readdata_21(ph_readdata_21),
	.ph_readdata_22(ph_readdata_22),
	.ph_readdata_23(ph_readdata_23),
	.ph_readdata_24(ph_readdata_24),
	.ph_readdata_25(ph_readdata_25),
	.ph_readdata_26(ph_readdata_26),
	.ph_readdata_27(ph_readdata_27),
	.ph_readdata_28(ph_readdata_28),
	.ph_readdata_29(ph_readdata_29),
	.ph_readdata_30(ph_readdata_30),
	.ph_readdata_31(ph_readdata_31),
	.mutex_grant(mutex_grant),
	.lif_waitrequest1(lif_waitrequest1),
	.lif_waitrequest2(lif_waitrequest2),
	.Equal8(Equal8),
	.basic_reconfig_waitrequest2(basic_reconfig_waitrequest2),
	.ctrl_go(ctrl_go),
	.ctrl_lock(ctrl_lock),
	.ctrl_opcode_2(ctrl_opcode_2),
	.ctrl_opcode_0(ctrl_opcode_0),
	.master_writedata_1(\inst_basic_acq|master_writedata[1]~q ),
	.master_writedata_2(\inst_basic_acq|master_writedata[2]~q ),
	.master_writedata_0(\inst_basic_acq|master_writedata[0]~q ),
	.master_writedata_3(\inst_basic_acq|master_writedata[3]~q ),
	.master_writedata_4(master_writedata_4),
	.master_writedata_5(master_writedata_5),
	.master_writedata_6(master_writedata_6),
	.master_writedata_7(master_writedata_7),
	.master_writedata_8(master_writedata_8),
	.master_writedata_9(master_writedata_9),
	.master_writedata_10(master_writedata_10),
	.master_writedata_11(master_writedata_11),
	.master_writedata_12(master_writedata_12),
	.master_writedata_13(master_writedata_13),
	.master_writedata_14(master_writedata_14),
	.master_writedata_15(master_writedata_15),
	.waitrequest_to_ctrl1(waitrequest_to_ctrl),
	.logical_ch_addr({ctrl_lch_9,ctrl_lch_8,ctrl_lch_7,ctrl_lch_6,ctrl_lch_5,ctrl_lch_4,ctrl_lch_3,ctrl_lch_2,ctrl_lch_1,ctrl_lch_0}),
	.ctrl_wdata_3(ctrl_wdata_3),
	.ctrl_wdata_4(ctrl_wdata_4),
	.ctrl_wdata_6(ctrl_wdata_6),
	.ctrl_wdata_7(ctrl_wdata_7),
	.ctrl_wdata_8(ctrl_wdata_8),
	.ctrl_wdata_10(ctrl_wdata_10),
	.ctrl_wdata_11(ctrl_wdata_11),
	.ctrl_wdata_12(ctrl_wdata_12),
	.readdata_for_user_0(readdata_for_user_0),
	.readdata_for_user_1(readdata_for_user_1),
	.readdata_for_user_2(readdata_for_user_2),
	.readdata_for_user_3(readdata_for_user_3),
	.readdata_for_user_4(readdata_for_user_4),
	.readdata_for_user_5(readdata_for_user_5),
	.readdata_for_user_6(readdata_for_user_6),
	.readdata_for_user_7(readdata_for_user_7),
	.readdata_for_user_8(readdata_for_user_8),
	.readdata_for_user_9(readdata_for_user_9),
	.readdata_for_user_10(readdata_for_user_10),
	.readdata_for_user_11(readdata_for_user_11),
	.readdata_for_user_12(readdata_for_user_12),
	.readdata_for_user_13(readdata_for_user_13),
	.readdata_for_user_14(readdata_for_user_14),
	.readdata_for_user_15(readdata_for_user_15),
	.readdata_for_user_16(readdata_for_user_16),
	.readdata_for_user_17(readdata_for_user_17),
	.readdata_for_user_18(readdata_for_user_18),
	.readdata_for_user_19(readdata_for_user_19),
	.readdata_for_user_20(readdata_for_user_20),
	.readdata_for_user_21(readdata_for_user_21),
	.readdata_for_user_22(readdata_for_user_22),
	.readdata_for_user_23(readdata_for_user_23),
	.readdata_for_user_24(readdata_for_user_24),
	.clk(mgmt_clk_clk));

endmodule

module RECONFIGURE_IP_alt_arbiter_acq_4 (
	grant_8,
	mutex_req,
	master_address_2,
	master_address_21,
	master_address_1,
	master_address_11,
	mutex_grant1,
	master_writedata_1,
	master_writedata_11,
	master_writedata_2,
	master_writedata_21,
	master_writedata_0,
	master_writedata_01,
	master_writedata_3,
	master_writedata_31)/* synthesis synthesis_greybox=0 */;
input 	grant_8;
input 	mutex_req;
input 	master_address_2;
output 	master_address_21;
input 	master_address_1;
output 	master_address_11;
output 	mutex_grant1;
input 	master_writedata_1;
output 	master_writedata_11;
input 	master_writedata_2;
output 	master_writedata_21;
input 	master_writedata_0;
output 	master_writedata_01;
input 	master_writedata_3;
output 	master_writedata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \master_address[2] (
	.dataa(!grant_8),
	.datab(!mutex_req),
	.datac(!master_address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_address_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_address[2] .extended_lut = "off";
defparam \master_address[2] .lut_mask = 64'h0101010101010101;
defparam \master_address[2] .shared_arith = "off";

cyclonev_lcell_comb \master_address[1] (
	.dataa(!grant_8),
	.datab(!mutex_req),
	.datac(!master_address_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_address_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_address[1] .extended_lut = "off";
defparam \master_address[1] .lut_mask = 64'h0101010101010101;
defparam \master_address[1] .shared_arith = "off";

cyclonev_lcell_comb mutex_grant(
	.dataa(!grant_8),
	.datab(!mutex_req),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mutex_grant1),
	.sumout(),
	.cout(),
	.shareout());
defparam mutex_grant.extended_lut = "off";
defparam mutex_grant.lut_mask = 64'h1111111111111111;
defparam mutex_grant.shared_arith = "off";

cyclonev_lcell_comb \master_writedata[1] (
	.dataa(!grant_8),
	.datab(!mutex_req),
	.datac(!master_writedata_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_writedata_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[1] .extended_lut = "off";
defparam \master_writedata[1] .lut_mask = 64'h0101010101010101;
defparam \master_writedata[1] .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[2] (
	.dataa(!grant_8),
	.datab(!mutex_req),
	.datac(!master_writedata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_writedata_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[2] .extended_lut = "off";
defparam \master_writedata[2] .lut_mask = 64'h0101010101010101;
defparam \master_writedata[2] .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[0] (
	.dataa(!grant_8),
	.datab(!mutex_req),
	.datac(!master_writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_writedata_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[0] .extended_lut = "off";
defparam \master_writedata[0] .lut_mask = 64'h0101010101010101;
defparam \master_writedata[0] .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[3] (
	.dataa(!grant_8),
	.datab(!mutex_req),
	.datac(!master_writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_writedata_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[3] .extended_lut = "off";
defparam \master_writedata[3] .lut_mask = 64'h0101010101010101;
defparam \master_writedata[3] .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_basic_acq_2 (
	basic_reconfig_readdata_12,
	basic_reconfig_readdata_13,
	basic_reconfig_readdata_14,
	basic_reconfig_readdata_15,
	basic_reconfig_readdata_16,
	basic_reconfig_readdata_17,
	basic_reconfig_readdata_18,
	basic_reconfig_readdata_19,
	basic_reconfig_readdata_20,
	basic_reconfig_readdata_21,
	basic_reconfig_readdata_22,
	basic_reconfig_readdata_23,
	basic_reconfig_readdata_24,
	basic_reconfig_readdata_25,
	basic_reconfig_readdata_26,
	basic_reconfig_readdata_27,
	basic_reconfig_readdata_28,
	basic_reconfig_readdata_29,
	basic_reconfig_readdata_30,
	basic_reconfig_readdata_31,
	ctrl_wdata_1,
	ctrl_addr_1,
	ctrl_wdata_2,
	ctrl_addr_5,
	ctrl_wdata_0,
	ctrl_addr_0,
	ctrl_addr_4,
	ctrl_wdata_5,
	ctrl_wdata_9,
	ctrl_wdata_13,
	ctrl_wdata_14,
	ctrl_wdata_15,
	basic_reconfig_readdata_0,
	basic_reconfig_readdata_1,
	basic_reconfig_readdata_2,
	basic_reconfig_readdata_3,
	basic_reconfig_readdata_4,
	basic_reconfig_readdata_5,
	basic_reconfig_readdata_6,
	basic_reconfig_readdata_7,
	basic_reconfig_readdata_8,
	basic_reconfig_readdata_9,
	basic_reconfig_readdata_10,
	basic_reconfig_readdata_11,
	master_write1,
	mutex_req1,
	master_address_2,
	master_address_0,
	master_address_1,
	lif_waitrequest,
	master_read1,
	basic_reconfig_waitrequest,
	basic_reconfig_waitrequest1,
	reset,
	ph_readdata_0,
	ph_readdata_1,
	ph_readdata_2,
	ph_readdata_3,
	ph_readdata_4,
	ph_readdata_5,
	ph_readdata_6,
	ph_readdata_7,
	ph_readdata_8,
	ph_readdata_9,
	illegal_phy_ch1,
	ph_readdata_10,
	ph_readdata_11,
	ph_readdata_12,
	ph_readdata_13,
	ph_readdata_14,
	ph_readdata_15,
	ph_readdata_16,
	ph_readdata_17,
	ph_readdata_18,
	ph_readdata_19,
	ph_readdata_20,
	ph_readdata_21,
	ph_readdata_22,
	ph_readdata_23,
	ph_readdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	mutex_grant,
	lif_waitrequest1,
	lif_waitrequest2,
	Equal8,
	basic_reconfig_waitrequest2,
	ctrl_go,
	ctrl_lock,
	ctrl_opcode_2,
	ctrl_opcode_0,
	master_writedata_1,
	master_writedata_2,
	master_writedata_0,
	master_writedata_3,
	master_writedata_4,
	master_writedata_5,
	master_writedata_6,
	master_writedata_7,
	master_writedata_8,
	master_writedata_9,
	master_writedata_10,
	master_writedata_11,
	master_writedata_12,
	master_writedata_13,
	master_writedata_14,
	master_writedata_15,
	waitrequest_to_ctrl1,
	logical_ch_addr,
	ctrl_wdata_3,
	ctrl_wdata_4,
	ctrl_wdata_6,
	ctrl_wdata_7,
	ctrl_wdata_8,
	ctrl_wdata_10,
	ctrl_wdata_11,
	ctrl_wdata_12,
	readdata_for_user_0,
	readdata_for_user_1,
	readdata_for_user_2,
	readdata_for_user_3,
	readdata_for_user_4,
	readdata_for_user_5,
	readdata_for_user_6,
	readdata_for_user_7,
	readdata_for_user_8,
	readdata_for_user_9,
	readdata_for_user_10,
	readdata_for_user_11,
	readdata_for_user_12,
	readdata_for_user_13,
	readdata_for_user_14,
	readdata_for_user_15,
	readdata_for_user_16,
	readdata_for_user_17,
	readdata_for_user_18,
	readdata_for_user_19,
	readdata_for_user_20,
	readdata_for_user_21,
	readdata_for_user_22,
	readdata_for_user_23,
	readdata_for_user_24,
	clk)/* synthesis synthesis_greybox=0 */;
input 	basic_reconfig_readdata_12;
input 	basic_reconfig_readdata_13;
input 	basic_reconfig_readdata_14;
input 	basic_reconfig_readdata_15;
input 	basic_reconfig_readdata_16;
input 	basic_reconfig_readdata_17;
input 	basic_reconfig_readdata_18;
input 	basic_reconfig_readdata_19;
input 	basic_reconfig_readdata_20;
input 	basic_reconfig_readdata_21;
input 	basic_reconfig_readdata_22;
input 	basic_reconfig_readdata_23;
input 	basic_reconfig_readdata_24;
input 	basic_reconfig_readdata_25;
input 	basic_reconfig_readdata_26;
input 	basic_reconfig_readdata_27;
input 	basic_reconfig_readdata_28;
input 	basic_reconfig_readdata_29;
input 	basic_reconfig_readdata_30;
input 	basic_reconfig_readdata_31;
input 	ctrl_wdata_1;
input 	ctrl_addr_1;
input 	ctrl_wdata_2;
input 	ctrl_addr_5;
input 	ctrl_wdata_0;
input 	ctrl_addr_0;
input 	ctrl_addr_4;
input 	ctrl_wdata_5;
input 	ctrl_wdata_9;
input 	ctrl_wdata_13;
input 	ctrl_wdata_14;
input 	ctrl_wdata_15;
input 	basic_reconfig_readdata_0;
input 	basic_reconfig_readdata_1;
input 	basic_reconfig_readdata_2;
input 	basic_reconfig_readdata_3;
input 	basic_reconfig_readdata_4;
input 	basic_reconfig_readdata_5;
input 	basic_reconfig_readdata_6;
input 	basic_reconfig_readdata_7;
input 	basic_reconfig_readdata_8;
input 	basic_reconfig_readdata_9;
input 	basic_reconfig_readdata_10;
input 	basic_reconfig_readdata_11;
output 	master_write1;
output 	mutex_req1;
output 	master_address_2;
output 	master_address_0;
output 	master_address_1;
input 	lif_waitrequest;
output 	master_read1;
input 	basic_reconfig_waitrequest;
input 	basic_reconfig_waitrequest1;
input 	reset;
output 	ph_readdata_0;
output 	ph_readdata_1;
output 	ph_readdata_2;
output 	ph_readdata_3;
output 	ph_readdata_4;
output 	ph_readdata_5;
output 	ph_readdata_6;
output 	ph_readdata_7;
output 	ph_readdata_8;
output 	ph_readdata_9;
output 	illegal_phy_ch1;
output 	ph_readdata_10;
output 	ph_readdata_11;
output 	ph_readdata_12;
output 	ph_readdata_13;
output 	ph_readdata_14;
output 	ph_readdata_15;
output 	ph_readdata_16;
output 	ph_readdata_17;
output 	ph_readdata_18;
output 	ph_readdata_19;
output 	ph_readdata_20;
output 	ph_readdata_21;
output 	ph_readdata_22;
output 	ph_readdata_23;
output 	ph_readdata_24;
output 	ph_readdata_25;
output 	ph_readdata_26;
output 	ph_readdata_27;
output 	ph_readdata_28;
output 	ph_readdata_29;
output 	ph_readdata_30;
output 	ph_readdata_31;
input 	mutex_grant;
input 	lif_waitrequest1;
input 	lif_waitrequest2;
output 	Equal8;
input 	basic_reconfig_waitrequest2;
input 	ctrl_go;
input 	ctrl_lock;
input 	ctrl_opcode_2;
input 	ctrl_opcode_0;
output 	master_writedata_1;
output 	master_writedata_2;
output 	master_writedata_0;
output 	master_writedata_3;
output 	master_writedata_4;
output 	master_writedata_5;
output 	master_writedata_6;
output 	master_writedata_7;
output 	master_writedata_8;
output 	master_writedata_9;
output 	master_writedata_10;
output 	master_writedata_11;
output 	master_writedata_12;
output 	master_writedata_13;
output 	master_writedata_14;
output 	master_writedata_15;
output 	waitrequest_to_ctrl1;
input 	[9:0] logical_ch_addr;
input 	ctrl_wdata_3;
input 	ctrl_wdata_4;
input 	ctrl_wdata_6;
input 	ctrl_wdata_7;
input 	ctrl_wdata_8;
input 	ctrl_wdata_10;
input 	ctrl_wdata_11;
input 	ctrl_wdata_12;
output 	readdata_for_user_0;
output 	readdata_for_user_1;
output 	readdata_for_user_2;
output 	readdata_for_user_3;
output 	readdata_for_user_4;
output 	readdata_for_user_5;
output 	readdata_for_user_6;
output 	readdata_for_user_7;
output 	readdata_for_user_8;
output 	readdata_for_user_9;
output 	readdata_for_user_10;
output 	readdata_for_user_11;
output 	readdata_for_user_12;
output 	readdata_for_user_13;
output 	readdata_for_user_14;
output 	readdata_for_user_15;
output 	readdata_for_user_16;
output 	readdata_for_user_17;
output 	readdata_for_user_18;
output 	readdata_for_user_19;
output 	readdata_for_user_20;
output 	readdata_for_user_21;
output 	readdata_for_user_22;
output 	readdata_for_user_23;
output 	readdata_for_user_24;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state.ST_READ_RECONFIG_BASIC_DATA~q ;
wire \lch_dly[4]~q ;
wire \lch_dly[5]~q ;
wire \lch_dly[2]~q ;
wire \lch_dly[3]~q ;
wire \lch_dly[0]~q ;
wire \lch_dly[1]~q ;
wire \lch_legal~0_combout ;
wire \lch_legal~1_combout ;
wire \lch_legal~2_combout ;
wire \lch_dly[8]~q ;
wire \lch_dly[9]~q ;
wire \lch_dly[6]~q ;
wire \lch_dly[7]~q ;
wire \lch_legal~3_combout ;
wire \lch_legal~4_combout ;
wire \lch_legal~5_combout ;
wire \lch_legal~q ;
wire \Selector3~5_combout ;
wire \master_writedata[5]~0_combout ;
wire \Selector8~0_combout ;
wire \Selector8~1_combout ;
wire \state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ;
wire \Selector9~0_combout ;
wire \state.ST_SET_RECONFIG_BASIC_WRITE~q ;
wire \phy_addr_is_set~0_combout ;
wire \phy_addr_is_set~q ;
wire \Selector3~9_combout ;
wire \Selector13~0_combout ;
wire \state.ST_START_AGAIN~q ;
wire \Selector15~0_combout ;
wire \Selector3~11_combout ;
wire \Selector3~13_combout ;
wire \Selector5~1_combout ;
wire \Selector5~2_combout ;
wire \state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ;
wire \Selector3~6_combout ;
wire \Selector3~8_combout ;
wire \Selector3~10_combout ;
wire \Selector15~1_combout ;
wire \Selector3~12_combout ;
wire \Selector15~2_combout ;
wire \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ;
wire \Selector12~0_combout ;
wire \Selector12~1_combout ;
wire \state.ST_CHECK_CTRLLOCK~q ;
wire \Selector14~0_combout ;
wire \state.ST_RELEASE_REQ~q ;
wire \Selector0~0_combout ;
wire \state.0000~q ;
wire \Selector1~0_combout ;
wire \state.ST_REQ_MUTEX~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \state.ST_WRITE_RECONFIG_BASIC_LCH~q ;
wire \Selector3~4_combout ;
wire \Selector3~7_combout ;
wire \state.ST_READ_PHY_ADDRESS~q ;
wire \Selector4~0_combout ;
wire \state.ST_CHECK_PHY_ADD_LEGAL~q ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ;
wire \Selector10~0_combout ;
wire \state.ST_SET_RECONFIG_BASIC_READ~q ;
wire \Selector11~0_combout ;
wire \WideOr17~0_combout ;
wire \WideOr7~0_combout ;
wire \WideOr8~combout ;
wire \Selector5~0_combout ;
wire \WideOr6~0_combout ;
wire \WideOr6~1_combout ;
wire \master_writedata[5]~1_combout ;
wire \WideOr5~0_combout ;
wire \WideOr17~1_combout ;
wire \Selector29~0_combout ;
wire \WideOr7~combout ;
wire \WideOr6~combout ;
wire \WideOr9~combout ;
wire \ph_readdata[13]~0_combout ;
wire \Selector16~0_combout ;
wire \ph_readdata[13]~1_combout ;
wire \Selector27~0_combout ;
wire \Selector27~1_combout ;
wire \Selector27~2_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \Selector28~0_combout ;
wire \Selector28~1_combout ;
wire \Selector25~0_combout ;
wire \master_writedata[5]~2_combout ;
wire \master_writedata[5]~3_combout ;
wire \Selector24~0_combout ;
wire \Selector23~0_combout ;
wire \Selector22~0_combout ;
wire \Selector21~0_combout ;
wire \Selector20~0_combout ;
wire \Selector19~0_combout ;
wire \Selector18~0_combout ;
wire \Selector17~0_combout ;
wire \master_writedata~4_combout ;
wire \master_writedata~5_combout ;
wire \master_writedata~6_combout ;
wire \master_writedata~7_combout ;
wire \Selector16~1_combout ;
wire \Selector16~2_combout ;
wire \readdata_for_user[0]~0_combout ;


dffeas master_write(
	.clk(clk),
	.d(\WideOr8~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_write1),
	.prn(vcc));
defparam master_write.is_wysiwyg = "true";
defparam master_write.power_up = "low";

dffeas mutex_req(
	.clk(clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mutex_req1),
	.prn(vcc));
defparam mutex_req.is_wysiwyg = "true";
defparam mutex_req.power_up = "low";

dffeas \master_address[2] (
	.clk(clk),
	.d(\WideOr5~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_2),
	.prn(vcc));
defparam \master_address[2] .is_wysiwyg = "true";
defparam \master_address[2] .power_up = "low";

dffeas \master_address[0] (
	.clk(clk),
	.d(\WideOr7~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_0),
	.prn(vcc));
defparam \master_address[0] .is_wysiwyg = "true";
defparam \master_address[0] .power_up = "low";

dffeas \master_address[1] (
	.clk(clk),
	.d(\WideOr6~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_address_1),
	.prn(vcc));
defparam \master_address[1] .is_wysiwyg = "true";
defparam \master_address[1] .power_up = "low";

dffeas master_read(
	.clk(clk),
	.d(\WideOr9~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_read1),
	.prn(vcc));
defparam master_read.is_wysiwyg = "true";
defparam master_read.power_up = "low";

dffeas \ph_readdata[0] (
	.clk(clk),
	.d(basic_reconfig_readdata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_0),
	.prn(vcc));
defparam \ph_readdata[0] .is_wysiwyg = "true";
defparam \ph_readdata[0] .power_up = "low";

dffeas \ph_readdata[1] (
	.clk(clk),
	.d(basic_reconfig_readdata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_1),
	.prn(vcc));
defparam \ph_readdata[1] .is_wysiwyg = "true";
defparam \ph_readdata[1] .power_up = "low";

dffeas \ph_readdata[2] (
	.clk(clk),
	.d(basic_reconfig_readdata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_2),
	.prn(vcc));
defparam \ph_readdata[2] .is_wysiwyg = "true";
defparam \ph_readdata[2] .power_up = "low";

dffeas \ph_readdata[3] (
	.clk(clk),
	.d(basic_reconfig_readdata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_3),
	.prn(vcc));
defparam \ph_readdata[3] .is_wysiwyg = "true";
defparam \ph_readdata[3] .power_up = "low";

dffeas \ph_readdata[4] (
	.clk(clk),
	.d(basic_reconfig_readdata_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_4),
	.prn(vcc));
defparam \ph_readdata[4] .is_wysiwyg = "true";
defparam \ph_readdata[4] .power_up = "low";

dffeas \ph_readdata[5] (
	.clk(clk),
	.d(basic_reconfig_readdata_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_5),
	.prn(vcc));
defparam \ph_readdata[5] .is_wysiwyg = "true";
defparam \ph_readdata[5] .power_up = "low";

dffeas \ph_readdata[6] (
	.clk(clk),
	.d(basic_reconfig_readdata_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_6),
	.prn(vcc));
defparam \ph_readdata[6] .is_wysiwyg = "true";
defparam \ph_readdata[6] .power_up = "low";

dffeas \ph_readdata[7] (
	.clk(clk),
	.d(basic_reconfig_readdata_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_7),
	.prn(vcc));
defparam \ph_readdata[7] .is_wysiwyg = "true";
defparam \ph_readdata[7] .power_up = "low";

dffeas \ph_readdata[8] (
	.clk(clk),
	.d(basic_reconfig_readdata_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_8),
	.prn(vcc));
defparam \ph_readdata[8] .is_wysiwyg = "true";
defparam \ph_readdata[8] .power_up = "low";

dffeas \ph_readdata[9] (
	.clk(clk),
	.d(basic_reconfig_readdata_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_9),
	.prn(vcc));
defparam \ph_readdata[9] .is_wysiwyg = "true";
defparam \ph_readdata[9] .power_up = "low";

dffeas illegal_phy_ch(
	.clk(clk),
	.d(Equal8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(illegal_phy_ch1),
	.prn(vcc));
defparam illegal_phy_ch.is_wysiwyg = "true";
defparam illegal_phy_ch.power_up = "low";

dffeas \ph_readdata[10] (
	.clk(clk),
	.d(basic_reconfig_readdata_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_10),
	.prn(vcc));
defparam \ph_readdata[10] .is_wysiwyg = "true";
defparam \ph_readdata[10] .power_up = "low";

dffeas \ph_readdata[11] (
	.clk(clk),
	.d(basic_reconfig_readdata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_11),
	.prn(vcc));
defparam \ph_readdata[11] .is_wysiwyg = "true";
defparam \ph_readdata[11] .power_up = "low";

dffeas \ph_readdata[12] (
	.clk(clk),
	.d(basic_reconfig_readdata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_12),
	.prn(vcc));
defparam \ph_readdata[12] .is_wysiwyg = "true";
defparam \ph_readdata[12] .power_up = "low";

dffeas \ph_readdata[13] (
	.clk(clk),
	.d(basic_reconfig_readdata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_13),
	.prn(vcc));
defparam \ph_readdata[13] .is_wysiwyg = "true";
defparam \ph_readdata[13] .power_up = "low";

dffeas \ph_readdata[14] (
	.clk(clk),
	.d(basic_reconfig_readdata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_14),
	.prn(vcc));
defparam \ph_readdata[14] .is_wysiwyg = "true";
defparam \ph_readdata[14] .power_up = "low";

dffeas \ph_readdata[15] (
	.clk(clk),
	.d(basic_reconfig_readdata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_15),
	.prn(vcc));
defparam \ph_readdata[15] .is_wysiwyg = "true";
defparam \ph_readdata[15] .power_up = "low";

dffeas \ph_readdata[16] (
	.clk(clk),
	.d(basic_reconfig_readdata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_16),
	.prn(vcc));
defparam \ph_readdata[16] .is_wysiwyg = "true";
defparam \ph_readdata[16] .power_up = "low";

dffeas \ph_readdata[17] (
	.clk(clk),
	.d(basic_reconfig_readdata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_17),
	.prn(vcc));
defparam \ph_readdata[17] .is_wysiwyg = "true";
defparam \ph_readdata[17] .power_up = "low";

dffeas \ph_readdata[18] (
	.clk(clk),
	.d(basic_reconfig_readdata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_18),
	.prn(vcc));
defparam \ph_readdata[18] .is_wysiwyg = "true";
defparam \ph_readdata[18] .power_up = "low";

dffeas \ph_readdata[19] (
	.clk(clk),
	.d(basic_reconfig_readdata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_19),
	.prn(vcc));
defparam \ph_readdata[19] .is_wysiwyg = "true";
defparam \ph_readdata[19] .power_up = "low";

dffeas \ph_readdata[20] (
	.clk(clk),
	.d(basic_reconfig_readdata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_20),
	.prn(vcc));
defparam \ph_readdata[20] .is_wysiwyg = "true";
defparam \ph_readdata[20] .power_up = "low";

dffeas \ph_readdata[21] (
	.clk(clk),
	.d(basic_reconfig_readdata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_21),
	.prn(vcc));
defparam \ph_readdata[21] .is_wysiwyg = "true";
defparam \ph_readdata[21] .power_up = "low";

dffeas \ph_readdata[22] (
	.clk(clk),
	.d(basic_reconfig_readdata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_22),
	.prn(vcc));
defparam \ph_readdata[22] .is_wysiwyg = "true";
defparam \ph_readdata[22] .power_up = "low";

dffeas \ph_readdata[23] (
	.clk(clk),
	.d(basic_reconfig_readdata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_23),
	.prn(vcc));
defparam \ph_readdata[23] .is_wysiwyg = "true";
defparam \ph_readdata[23] .power_up = "low";

dffeas \ph_readdata[24] (
	.clk(clk),
	.d(basic_reconfig_readdata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_24),
	.prn(vcc));
defparam \ph_readdata[24] .is_wysiwyg = "true";
defparam \ph_readdata[24] .power_up = "low";

dffeas \ph_readdata[25] (
	.clk(clk),
	.d(basic_reconfig_readdata_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_25),
	.prn(vcc));
defparam \ph_readdata[25] .is_wysiwyg = "true";
defparam \ph_readdata[25] .power_up = "low";

dffeas \ph_readdata[26] (
	.clk(clk),
	.d(basic_reconfig_readdata_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_26),
	.prn(vcc));
defparam \ph_readdata[26] .is_wysiwyg = "true";
defparam \ph_readdata[26] .power_up = "low";

dffeas \ph_readdata[27] (
	.clk(clk),
	.d(basic_reconfig_readdata_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_27),
	.prn(vcc));
defparam \ph_readdata[27] .is_wysiwyg = "true";
defparam \ph_readdata[27] .power_up = "low";

dffeas \ph_readdata[28] (
	.clk(clk),
	.d(basic_reconfig_readdata_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_28),
	.prn(vcc));
defparam \ph_readdata[28] .is_wysiwyg = "true";
defparam \ph_readdata[28] .power_up = "low";

dffeas \ph_readdata[29] (
	.clk(clk),
	.d(basic_reconfig_readdata_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_29),
	.prn(vcc));
defparam \ph_readdata[29] .is_wysiwyg = "true";
defparam \ph_readdata[29] .power_up = "low";

dffeas \ph_readdata[30] (
	.clk(clk),
	.d(basic_reconfig_readdata_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_30),
	.prn(vcc));
defparam \ph_readdata[30] .is_wysiwyg = "true";
defparam \ph_readdata[30] .power_up = "low";

dffeas \ph_readdata[31] (
	.clk(clk),
	.d(basic_reconfig_readdata_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ph_readdata[13]~1_combout ),
	.q(ph_readdata_31),
	.prn(vcc));
defparam \ph_readdata[31] .is_wysiwyg = "true";
defparam \ph_readdata[31] .power_up = "low";

cyclonev_lcell_comb \Equal8~0 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!basic_reconfig_readdata_1),
	.datac(!basic_reconfig_readdata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal8),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal8~0 .extended_lut = "off";
defparam \Equal8~0 .lut_mask = 64'h0101010101010101;
defparam \Equal8~0 .shared_arith = "off";

dffeas \master_writedata[1] (
	.clk(clk),
	.d(\Selector27~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_1),
	.prn(vcc));
defparam \master_writedata[1] .is_wysiwyg = "true";
defparam \master_writedata[1] .power_up = "low";

dffeas \master_writedata[2] (
	.clk(clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_2),
	.prn(vcc));
defparam \master_writedata[2] .is_wysiwyg = "true";
defparam \master_writedata[2] .power_up = "low";

dffeas \master_writedata[0] (
	.clk(clk),
	.d(\Selector28~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_0),
	.prn(vcc));
defparam \master_writedata[0] .is_wysiwyg = "true";
defparam \master_writedata[0] .power_up = "low";

dffeas \master_writedata[3] (
	.clk(clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_3),
	.prn(vcc));
defparam \master_writedata[3] .is_wysiwyg = "true";
defparam \master_writedata[3] .power_up = "low";

dffeas \master_writedata[4] (
	.clk(clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_4),
	.prn(vcc));
defparam \master_writedata[4] .is_wysiwyg = "true";
defparam \master_writedata[4] .power_up = "low";

dffeas \master_writedata[5] (
	.clk(clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_5),
	.prn(vcc));
defparam \master_writedata[5] .is_wysiwyg = "true";
defparam \master_writedata[5] .power_up = "low";

dffeas \master_writedata[6] (
	.clk(clk),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_6),
	.prn(vcc));
defparam \master_writedata[6] .is_wysiwyg = "true";
defparam \master_writedata[6] .power_up = "low";

dffeas \master_writedata[7] (
	.clk(clk),
	.d(\Selector21~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_7),
	.prn(vcc));
defparam \master_writedata[7] .is_wysiwyg = "true";
defparam \master_writedata[7] .power_up = "low";

dffeas \master_writedata[8] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_8),
	.prn(vcc));
defparam \master_writedata[8] .is_wysiwyg = "true";
defparam \master_writedata[8] .power_up = "low";

dffeas \master_writedata[9] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_9),
	.prn(vcc));
defparam \master_writedata[9] .is_wysiwyg = "true";
defparam \master_writedata[9] .power_up = "low";

dffeas \master_writedata[10] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_10),
	.prn(vcc));
defparam \master_writedata[10] .is_wysiwyg = "true";
defparam \master_writedata[10] .power_up = "low";

dffeas \master_writedata[11] (
	.clk(clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_11),
	.prn(vcc));
defparam \master_writedata[11] .is_wysiwyg = "true";
defparam \master_writedata[11] .power_up = "low";

dffeas \master_writedata[12] (
	.clk(clk),
	.d(\master_writedata~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_12),
	.prn(vcc));
defparam \master_writedata[12] .is_wysiwyg = "true";
defparam \master_writedata[12] .power_up = "low";

dffeas \master_writedata[13] (
	.clk(clk),
	.d(\master_writedata~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_13),
	.prn(vcc));
defparam \master_writedata[13] .is_wysiwyg = "true";
defparam \master_writedata[13] .power_up = "low";

dffeas \master_writedata[14] (
	.clk(clk),
	.d(\master_writedata~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_14),
	.prn(vcc));
defparam \master_writedata[14] .is_wysiwyg = "true";
defparam \master_writedata[14] .power_up = "low";

dffeas \master_writedata[15] (
	.clk(clk),
	.d(\master_writedata~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(master_writedata_15),
	.prn(vcc));
defparam \master_writedata[15] .is_wysiwyg = "true";
defparam \master_writedata[15] .power_up = "low";

dffeas waitrequest_to_ctrl(
	.clk(clk),
	.d(\Selector16~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_to_ctrl1),
	.prn(vcc));
defparam waitrequest_to_ctrl.is_wysiwyg = "true";
defparam waitrequest_to_ctrl.power_up = "low";

dffeas \readdata_for_user[0] (
	.clk(clk),
	.d(basic_reconfig_readdata_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_0),
	.prn(vcc));
defparam \readdata_for_user[0] .is_wysiwyg = "true";
defparam \readdata_for_user[0] .power_up = "low";

dffeas \readdata_for_user[1] (
	.clk(clk),
	.d(basic_reconfig_readdata_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_1),
	.prn(vcc));
defparam \readdata_for_user[1] .is_wysiwyg = "true";
defparam \readdata_for_user[1] .power_up = "low";

dffeas \readdata_for_user[2] (
	.clk(clk),
	.d(basic_reconfig_readdata_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_2),
	.prn(vcc));
defparam \readdata_for_user[2] .is_wysiwyg = "true";
defparam \readdata_for_user[2] .power_up = "low";

dffeas \readdata_for_user[3] (
	.clk(clk),
	.d(basic_reconfig_readdata_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_3),
	.prn(vcc));
defparam \readdata_for_user[3] .is_wysiwyg = "true";
defparam \readdata_for_user[3] .power_up = "low";

dffeas \readdata_for_user[4] (
	.clk(clk),
	.d(basic_reconfig_readdata_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_4),
	.prn(vcc));
defparam \readdata_for_user[4] .is_wysiwyg = "true";
defparam \readdata_for_user[4] .power_up = "low";

dffeas \readdata_for_user[5] (
	.clk(clk),
	.d(basic_reconfig_readdata_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_5),
	.prn(vcc));
defparam \readdata_for_user[5] .is_wysiwyg = "true";
defparam \readdata_for_user[5] .power_up = "low";

dffeas \readdata_for_user[6] (
	.clk(clk),
	.d(basic_reconfig_readdata_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_6),
	.prn(vcc));
defparam \readdata_for_user[6] .is_wysiwyg = "true";
defparam \readdata_for_user[6] .power_up = "low";

dffeas \readdata_for_user[7] (
	.clk(clk),
	.d(basic_reconfig_readdata_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_7),
	.prn(vcc));
defparam \readdata_for_user[7] .is_wysiwyg = "true";
defparam \readdata_for_user[7] .power_up = "low";

dffeas \readdata_for_user[8] (
	.clk(clk),
	.d(basic_reconfig_readdata_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_8),
	.prn(vcc));
defparam \readdata_for_user[8] .is_wysiwyg = "true";
defparam \readdata_for_user[8] .power_up = "low";

dffeas \readdata_for_user[9] (
	.clk(clk),
	.d(basic_reconfig_readdata_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_9),
	.prn(vcc));
defparam \readdata_for_user[9] .is_wysiwyg = "true";
defparam \readdata_for_user[9] .power_up = "low";

dffeas \readdata_for_user[10] (
	.clk(clk),
	.d(basic_reconfig_readdata_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_10),
	.prn(vcc));
defparam \readdata_for_user[10] .is_wysiwyg = "true";
defparam \readdata_for_user[10] .power_up = "low";

dffeas \readdata_for_user[11] (
	.clk(clk),
	.d(basic_reconfig_readdata_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_11),
	.prn(vcc));
defparam \readdata_for_user[11] .is_wysiwyg = "true";
defparam \readdata_for_user[11] .power_up = "low";

dffeas \readdata_for_user[12] (
	.clk(clk),
	.d(basic_reconfig_readdata_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_12),
	.prn(vcc));
defparam \readdata_for_user[12] .is_wysiwyg = "true";
defparam \readdata_for_user[12] .power_up = "low";

dffeas \readdata_for_user[13] (
	.clk(clk),
	.d(basic_reconfig_readdata_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_13),
	.prn(vcc));
defparam \readdata_for_user[13] .is_wysiwyg = "true";
defparam \readdata_for_user[13] .power_up = "low";

dffeas \readdata_for_user[14] (
	.clk(clk),
	.d(basic_reconfig_readdata_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_14),
	.prn(vcc));
defparam \readdata_for_user[14] .is_wysiwyg = "true";
defparam \readdata_for_user[14] .power_up = "low";

dffeas \readdata_for_user[15] (
	.clk(clk),
	.d(basic_reconfig_readdata_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_15),
	.prn(vcc));
defparam \readdata_for_user[15] .is_wysiwyg = "true";
defparam \readdata_for_user[15] .power_up = "low";

dffeas \readdata_for_user[16] (
	.clk(clk),
	.d(basic_reconfig_readdata_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_16),
	.prn(vcc));
defparam \readdata_for_user[16] .is_wysiwyg = "true";
defparam \readdata_for_user[16] .power_up = "low";

dffeas \readdata_for_user[17] (
	.clk(clk),
	.d(basic_reconfig_readdata_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_17),
	.prn(vcc));
defparam \readdata_for_user[17] .is_wysiwyg = "true";
defparam \readdata_for_user[17] .power_up = "low";

dffeas \readdata_for_user[18] (
	.clk(clk),
	.d(basic_reconfig_readdata_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_18),
	.prn(vcc));
defparam \readdata_for_user[18] .is_wysiwyg = "true";
defparam \readdata_for_user[18] .power_up = "low";

dffeas \readdata_for_user[19] (
	.clk(clk),
	.d(basic_reconfig_readdata_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_19),
	.prn(vcc));
defparam \readdata_for_user[19] .is_wysiwyg = "true";
defparam \readdata_for_user[19] .power_up = "low";

dffeas \readdata_for_user[20] (
	.clk(clk),
	.d(basic_reconfig_readdata_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_20),
	.prn(vcc));
defparam \readdata_for_user[20] .is_wysiwyg = "true";
defparam \readdata_for_user[20] .power_up = "low";

dffeas \readdata_for_user[21] (
	.clk(clk),
	.d(basic_reconfig_readdata_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_21),
	.prn(vcc));
defparam \readdata_for_user[21] .is_wysiwyg = "true";
defparam \readdata_for_user[21] .power_up = "low";

dffeas \readdata_for_user[22] (
	.clk(clk),
	.d(basic_reconfig_readdata_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_22),
	.prn(vcc));
defparam \readdata_for_user[22] .is_wysiwyg = "true";
defparam \readdata_for_user[22] .power_up = "low";

dffeas \readdata_for_user[23] (
	.clk(clk),
	.d(basic_reconfig_readdata_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_23),
	.prn(vcc));
defparam \readdata_for_user[23] .is_wysiwyg = "true";
defparam \readdata_for_user[23] .power_up = "low";

dffeas \readdata_for_user[24] (
	.clk(clk),
	.d(basic_reconfig_readdata_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_for_user[0]~0_combout ),
	.q(readdata_for_user_24),
	.prn(vcc));
defparam \readdata_for_user[24] .is_wysiwyg = "true";
defparam \readdata_for_user[24] .power_up = "low";

dffeas \state.ST_READ_RECONFIG_BASIC_DATA (
	.clk(clk),
	.d(\Selector11~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.prn(vcc));
defparam \state.ST_READ_RECONFIG_BASIC_DATA .is_wysiwyg = "true";
defparam \state.ST_READ_RECONFIG_BASIC_DATA .power_up = "low";

dffeas \lch_dly[4] (
	.clk(clk),
	.d(logical_ch_addr[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[4]~q ),
	.prn(vcc));
defparam \lch_dly[4] .is_wysiwyg = "true";
defparam \lch_dly[4] .power_up = "low";

dffeas \lch_dly[5] (
	.clk(clk),
	.d(logical_ch_addr[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[5]~q ),
	.prn(vcc));
defparam \lch_dly[5] .is_wysiwyg = "true";
defparam \lch_dly[5] .power_up = "low";

dffeas \lch_dly[2] (
	.clk(clk),
	.d(logical_ch_addr[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[2]~q ),
	.prn(vcc));
defparam \lch_dly[2] .is_wysiwyg = "true";
defparam \lch_dly[2] .power_up = "low";

dffeas \lch_dly[3] (
	.clk(clk),
	.d(logical_ch_addr[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[3]~q ),
	.prn(vcc));
defparam \lch_dly[3] .is_wysiwyg = "true";
defparam \lch_dly[3] .power_up = "low";

dffeas \lch_dly[0] (
	.clk(clk),
	.d(logical_ch_addr[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[0]~q ),
	.prn(vcc));
defparam \lch_dly[0] .is_wysiwyg = "true";
defparam \lch_dly[0] .power_up = "low";

dffeas \lch_dly[1] (
	.clk(clk),
	.d(logical_ch_addr[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[1]~q ),
	.prn(vcc));
defparam \lch_dly[1] .is_wysiwyg = "true";
defparam \lch_dly[1] .power_up = "low";

cyclonev_lcell_comb \lch_legal~0 (
	.dataa(!\lch_dly[0]~q ),
	.datab(!logical_ch_addr[0]),
	.datac(!\lch_dly[1]~q ),
	.datad(!logical_ch_addr[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~0 .extended_lut = "off";
defparam \lch_legal~0 .lut_mask = 64'h9009900990099009;
defparam \lch_legal~0 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~1 (
	.dataa(!\lch_dly[2]~q ),
	.datab(!logical_ch_addr[2]),
	.datac(!\lch_dly[3]~q ),
	.datad(!logical_ch_addr[3]),
	.datae(!\lch_legal~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~1 .extended_lut = "off";
defparam \lch_legal~1 .lut_mask = 64'h0000900900009009;
defparam \lch_legal~1 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~2 (
	.dataa(!\lch_dly[4]~q ),
	.datab(!logical_ch_addr[4]),
	.datac(!\lch_dly[5]~q ),
	.datad(!logical_ch_addr[5]),
	.datae(!\lch_legal~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~2 .extended_lut = "off";
defparam \lch_legal~2 .lut_mask = 64'h0000900900009009;
defparam \lch_legal~2 .shared_arith = "off";

dffeas \lch_dly[8] (
	.clk(clk),
	.d(logical_ch_addr[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[8]~q ),
	.prn(vcc));
defparam \lch_dly[8] .is_wysiwyg = "true";
defparam \lch_dly[8] .power_up = "low";

dffeas \lch_dly[9] (
	.clk(clk),
	.d(logical_ch_addr[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[9]~q ),
	.prn(vcc));
defparam \lch_dly[9] .is_wysiwyg = "true";
defparam \lch_dly[9] .power_up = "low";

dffeas \lch_dly[6] (
	.clk(clk),
	.d(logical_ch_addr[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[6]~q ),
	.prn(vcc));
defparam \lch_dly[6] .is_wysiwyg = "true";
defparam \lch_dly[6] .power_up = "low";

dffeas \lch_dly[7] (
	.clk(clk),
	.d(logical_ch_addr[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_dly[7]~q ),
	.prn(vcc));
defparam \lch_dly[7] .is_wysiwyg = "true";
defparam \lch_dly[7] .power_up = "low";

cyclonev_lcell_comb \lch_legal~3 (
	.dataa(!\lch_dly[6]~q ),
	.datab(!logical_ch_addr[6]),
	.datac(!\lch_dly[7]~q ),
	.datad(!logical_ch_addr[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~3 .extended_lut = "off";
defparam \lch_legal~3 .lut_mask = 64'h9009900990099009;
defparam \lch_legal~3 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~4 (
	.dataa(!\lch_dly[8]~q ),
	.datab(!logical_ch_addr[8]),
	.datac(!\lch_dly[9]~q ),
	.datad(!logical_ch_addr[9]),
	.datae(!\lch_legal~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~4 .extended_lut = "off";
defparam \lch_legal~4 .lut_mask = 64'h0000900900009009;
defparam \lch_legal~4 .shared_arith = "off";

cyclonev_lcell_comb \lch_legal~5 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!Equal8),
	.datac(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datad(!\lch_legal~q ),
	.datae(!\lch_legal~2_combout ),
	.dataf(!\lch_legal~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lch_legal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lch_legal~5 .extended_lut = "off";
defparam \lch_legal~5 .lut_mask = 64'h00000000000008FF;
defparam \lch_legal~5 .shared_arith = "off";

dffeas lch_legal(
	.clk(clk),
	.d(\lch_legal~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\lch_legal~q ),
	.prn(vcc));
defparam lch_legal.is_wysiwyg = "true";
defparam lch_legal.power_up = "low";

cyclonev_lcell_comb \Selector3~5 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!basic_reconfig_readdata_1),
	.datac(!basic_reconfig_readdata_2),
	.datad(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~5 .extended_lut = "off";
defparam \Selector3~5 .lut_mask = 64'h0001000100010001;
defparam \Selector3~5 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[5]~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~5_combout ),
	.dataf(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[5]~0 .extended_lut = "off";
defparam \master_writedata[5]~0 .lut_mask = 64'hFFFF00007FFF0000;
defparam \master_writedata[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!ctrl_opcode_2),
	.datad(!ctrl_opcode_0),
	.datae(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h0000002000000020;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~1 (
	.dataa(!\master_writedata[5]~0_combout ),
	.datab(!\Selector3~8_combout ),
	.datac(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datad(!\Selector3~13_combout ),
	.datae(!\Selector8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~1 .extended_lut = "off";
defparam \Selector8~1 .lut_mask = 64'h0004FFBF0004FFBF;
defparam \Selector8~1 .shared_arith = "off";

dffeas \state.ST_WRITE_DATA_TO_RECONFIG_BASIC (
	.clk(clk),
	.d(\Selector8~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.prn(vcc));
defparam \state.ST_WRITE_DATA_TO_RECONFIG_BASIC .is_wysiwyg = "true";
defparam \state.ST_WRITE_DATA_TO_RECONFIG_BASIC .power_up = "low";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.dataf(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h00007FFF8000FFFF;
defparam \Selector9~0 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_WRITE (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_WRITE .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_WRITE .power_up = "low";

cyclonev_lcell_comb \phy_addr_is_set~0 (
	.dataa(!\phy_addr_is_set~q ),
	.datab(!\Selector15~2_combout ),
	.datac(!\Selector5~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\phy_addr_is_set~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \phy_addr_is_set~0 .extended_lut = "off";
defparam \phy_addr_is_set~0 .lut_mask = 64'h4C4C4C4C4C4C4C4C;
defparam \phy_addr_is_set~0 .shared_arith = "off";

dffeas phy_addr_is_set(
	.clk(clk),
	.d(\phy_addr_is_set~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\phy_addr_is_set~q ),
	.prn(vcc));
defparam phy_addr_is_set.is_wysiwyg = "true";
defparam phy_addr_is_set.power_up = "low";

cyclonev_lcell_comb \Selector3~9 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.datab(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.datac(!\phy_addr_is_set~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~9 .extended_lut = "off";
defparam \Selector3~9 .lut_mask = 64'h0707070707070707;
defparam \Selector3~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector13~0 (
	.dataa(!ctrl_go),
	.datab(!\state.ST_START_AGAIN~q ),
	.datac(!ctrl_lock),
	.datad(!\state.ST_CHECK_CTRLLOCK~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~0 .extended_lut = "off";
defparam \Selector13~0 .lut_mask = 64'h222F222F222F222F;
defparam \Selector13~0 .shared_arith = "off";

dffeas \state.ST_START_AGAIN (
	.clk(clk),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_START_AGAIN~q ),
	.prn(vcc));
defparam \state.ST_START_AGAIN .is_wysiwyg = "true";
defparam \state.ST_START_AGAIN .power_up = "low";

cyclonev_lcell_comb \Selector15~0 (
	.dataa(!\state.0000~q ),
	.datab(!\state.ST_REQ_MUTEX~q ),
	.datac(!\state.ST_START_AGAIN~q ),
	.datad(!\state.ST_CHECK_CTRLLOCK~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "off";
defparam \Selector15~0 .lut_mask = 64'h4000400040004000;
defparam \Selector15~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~11 (
	.dataa(!\Selector3~5_combout ),
	.datab(!\Selector3~4_combout ),
	.datac(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.datad(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~11 .extended_lut = "off";
defparam \Selector3~11 .lut_mask = 64'h8000800080008000;
defparam \Selector3~11 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~13 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\Selector3~4_combout ),
	.datad(!\Selector3~9_combout ),
	.datae(!\Selector15~0_combout ),
	.dataf(!\Selector3~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~13 .extended_lut = "off";
defparam \Selector3~13 .lut_mask = 64'h0000FDDD0000DDDD;
defparam \Selector3~13 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!ctrl_opcode_2),
	.datad(!ctrl_opcode_0),
	.datae(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'h0000000200000002;
defparam \Selector5~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~2 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.datab(!\master_writedata[5]~0_combout ),
	.datac(!\Selector3~8_combout ),
	.datad(!\Selector3~13_combout ),
	.datae(!\Selector5~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~2 .extended_lut = "off";
defparam \Selector5~2 .lut_mask = 64'h0010FFFF0010FFFF;
defparam \Selector5~2 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_PADDR_MODE (
	.clk(clk),
	.d(\Selector5~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_PADDR_MODE .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_PADDR_MODE .power_up = "low";

cyclonev_lcell_comb \Selector3~6 (
	.dataa(!ctrl_opcode_2),
	.datab(!ctrl_opcode_0),
	.datac(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~6 .extended_lut = "off";
defparam \Selector3~6 .lut_mask = 64'h0101010101010101;
defparam \Selector3~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~8 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~8 .extended_lut = "off";
defparam \Selector3~8 .lut_mask = 64'h0000800000008000;
defparam \Selector3~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~10 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~10 .extended_lut = "off";
defparam \Selector3~10 .lut_mask = 64'h0000800000008000;
defparam \Selector3~10 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~1 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~4_combout ),
	.dataf(!\Selector15~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~1 .extended_lut = "off";
defparam \Selector15~1 .lut_mask = 64'h00000000FFFF7FFF;
defparam \Selector15~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~12 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\Selector3~9_combout ),
	.dataf(!\Selector3~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~12 .extended_lut = "off";
defparam \Selector3~12 .lut_mask = 64'h0000000080000000;
defparam \Selector3~12 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~2 (
	.dataa(!\master_writedata[5]~0_combout ),
	.datab(!\Selector3~8_combout ),
	.datac(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datad(!\Selector3~10_combout ),
	.datae(!\Selector15~1_combout ),
	.dataf(!\Selector3~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~2 .extended_lut = "off";
defparam \Selector15~2 .lut_mask = 64'h0000044400000000;
defparam \Selector15~2 .shared_arith = "off";

dffeas \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE (
	.clk(clk),
	.d(\Selector15~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.prn(vcc));
defparam \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE .is_wysiwyg = "true";
defparam \state.ST_CLR_RECONFIG_BASIC_PADDR_MODE .power_up = "low";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_WRITE~q ),
	.datab(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'h8888888888888888;
defparam \Selector12~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~1 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_CHECK_CTRLLOCK~q ),
	.datad(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datae(!\Selector12~0_combout ),
	.dataf(!\phy_addr_is_set~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~1 .extended_lut = "off";
defparam \Selector12~1 .lut_mask = 64'h2F2F00220D2F0022;
defparam \Selector12~1 .shared_arith = "off";

dffeas \state.ST_CHECK_CTRLLOCK (
	.clk(clk),
	.d(\Selector12~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CHECK_CTRLLOCK~q ),
	.prn(vcc));
defparam \state.ST_CHECK_CTRLLOCK .is_wysiwyg = "true";
defparam \state.ST_CHECK_CTRLLOCK .power_up = "low";

cyclonev_lcell_comb \Selector14~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_RELEASE_REQ~q ),
	.datad(!ctrl_lock),
	.datae(!\state.ST_CHECK_CTRLLOCK~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~0 .extended_lut = "off";
defparam \Selector14~0 .lut_mask = 64'h0D0DFF0D0D0DFF0D;
defparam \Selector14~0 .shared_arith = "off";

dffeas \state.ST_RELEASE_REQ (
	.clk(clk),
	.d(\Selector14~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_RELEASE_REQ~q ),
	.prn(vcc));
defparam \state.ST_RELEASE_REQ .is_wysiwyg = "true";
defparam \state.ST_RELEASE_REQ .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_RELEASE_REQ~q ),
	.datad(!\Selector3~5_combout ),
	.datae(!ctrl_go),
	.dataf(!\state.0000~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h0000FD00FD00FD00;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.0000 (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.0000~q ),
	.prn(vcc));
defparam \state.0000 .is_wysiwyg = "true";
defparam \state.0000 .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!mutex_grant),
	.datab(!ctrl_go),
	.datac(!\state.0000~q ),
	.datad(!\state.ST_REQ_MUTEX~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h30BA30BA30BA30BA;
defparam \Selector1~0 .shared_arith = "off";

dffeas \state.ST_REQ_MUTEX (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_REQ_MUTEX~q ),
	.prn(vcc));
defparam \state.ST_REQ_MUTEX .is_wysiwyg = "true";
defparam \state.ST_REQ_MUTEX .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!mutex_grant),
	.datab(!\state.ST_REQ_MUTEX~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h1111111111111111;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h00007FFFFFFFFFFF;
defparam \Selector2~1 .shared_arith = "off";

dffeas \state.ST_WRITE_RECONFIG_BASIC_LCH (
	.clk(clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.prn(vcc));
defparam \state.ST_WRITE_RECONFIG_BASIC_LCH .is_wysiwyg = "true";
defparam \state.ST_WRITE_RECONFIG_BASIC_LCH .power_up = "low";

cyclonev_lcell_comb \Selector3~4 (
	.dataa(!\lch_legal~q ),
	.datab(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~4 .extended_lut = "off";
defparam \Selector3~4 .lut_mask = 64'h2222222222222222;
defparam \Selector3~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~7 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\Selector3~4_combout ),
	.datac(!\state.ST_READ_PHY_ADDRESS~q ),
	.datad(!\master_writedata[5]~0_combout ),
	.datae(!\Selector3~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~7 .extended_lut = "off";
defparam \Selector3~7 .lut_mask = 64'h0027000500270005;
defparam \Selector3~7 .shared_arith = "off";

dffeas \state.ST_READ_PHY_ADDRESS (
	.clk(clk),
	.d(\Selector3~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_READ_PHY_ADDRESS~q ),
	.prn(vcc));
defparam \state.ST_READ_PHY_ADDRESS .is_wysiwyg = "true";
defparam \state.ST_READ_PHY_ADDRESS .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!Equal8),
	.datac(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datad(!\state.ST_READ_PHY_ADDRESS~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h04AE04AE04AE04AE;
defparam \Selector4~0 .shared_arith = "off";

dffeas \state.ST_CHECK_PHY_ADD_LEGAL (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.prn(vcc));
defparam \state.ST_CHECK_PHY_ADD_LEGAL .is_wysiwyg = "true";
defparam \state.ST_CHECK_PHY_ADD_LEGAL .power_up = "low";

cyclonev_lcell_comb \Selector6~1 (
	.dataa(!Equal8),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!\lch_legal~q ),
	.datad(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'h222F222F222F222F;
defparam \Selector6~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~2 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.datae(!\Selector6~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~2 .extended_lut = "off";
defparam \Selector6~2 .lut_mask = 64'h00FB0CFF00FB0CFF;
defparam \Selector6~2 .shared_arith = "off";

dffeas \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK (
	.clk(clk),
	.d(\Selector6~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.prn(vcc));
defparam \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK .is_wysiwyg = "true";
defparam \state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK .power_up = "low";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!ctrl_go),
	.datab(!\state.ST_START_AGAIN~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h1111111111111111;
defparam \Selector7~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~1 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest1),
	.datad(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datae(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.dataf(!\Selector7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~1 .extended_lut = "off";
defparam \Selector7~1 .lut_mask = 64'h00F304F7FFFFFFFF;
defparam \Selector7~1 .shared_arith = "off";

dffeas \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG (
	.clk(clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.prn(vcc));
defparam \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG .is_wysiwyg = "true";
defparam \state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG .power_up = "low";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!ctrl_opcode_0),
	.datad(!\state.ST_ACCESS_RECONFIG_BASIC_OFFSET_REG~q ),
	.datae(!\Selector3~6_combout ),
	.dataf(!\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h00202222DDFDFFFF;
defparam \Selector10~0 .shared_arith = "off";

dffeas \state.ST_SET_RECONFIG_BASIC_READ (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.prn(vcc));
defparam \state.ST_SET_RECONFIG_BASIC_READ .is_wysiwyg = "true";
defparam \state.ST_SET_RECONFIG_BASIC_READ .power_up = "low";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!lif_waitrequest1),
	.datab(!lif_waitrequest),
	.datac(!basic_reconfig_waitrequest),
	.datad(!lif_waitrequest2),
	.datae(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.dataf(!\state.ST_SET_RECONFIG_BASIC_READ~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h00007FFF8000FFFF;
defparam \Selector11~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr17~0 (
	.dataa(!\Selector4~0_combout ),
	.datab(!\Selector12~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~0 .extended_lut = "off";
defparam \WideOr17~0 .lut_mask = 64'h8888888888888888;
defparam \WideOr17~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr7~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\Selector13~0_combout ),
	.datac(!\Selector3~7_combout ),
	.datad(!\WideOr17~0_combout ),
	.datae(!\Selector0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr7~0 .extended_lut = "off";
defparam \WideOr7~0 .lut_mask = 64'h0000008000000080;
defparam \WideOr7~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr8(
	.dataa(!\Selector11~0_combout ),
	.datab(!\Selector6~2_combout ),
	.datac(!\WideOr7~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr8~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr8.extended_lut = "off";
defparam WideOr8.lut_mask = 64'h0808080808080808;
defparam WideOr8.shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!\state.ST_SET_RECONFIG_BASIC_PADDR_MODE~q ),
	.datab(!\master_writedata[5]~0_combout ),
	.datac(!\Selector3~8_combout ),
	.datad(!\Selector3~10_combout ),
	.datae(!\Selector15~1_combout ),
	.dataf(!\Selector3~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h0000100000000000;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr6~0 (
	.dataa(!basic_reconfig_readdata_0),
	.datab(!basic_reconfig_waitrequest2),
	.datac(!\state.ST_CONFIRM_RECONFIG_BASIC_CH_LOCK~q ),
	.datad(!\Selector6~1_combout ),
	.datae(!\Selector9~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr6~0 .extended_lut = "off";
defparam \WideOr6~0 .lut_mask = 64'hF4300000F4300000;
defparam \WideOr6~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr6~1 (
	.dataa(!\Selector3~7_combout ),
	.datab(!\Selector15~2_combout ),
	.datac(!\Selector5~0_combout ),
	.datad(!\Selector5~1_combout ),
	.datae(!\Selector10~0_combout ),
	.dataf(!\WideOr6~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr6~1 .extended_lut = "off";
defparam \WideOr6~1 .lut_mask = 64'h0000000080000000;
defparam \WideOr6~1 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[5]~1 (
	.dataa(!\master_writedata[5]~0_combout ),
	.datab(!\Selector3~10_combout ),
	.datac(!\Selector15~1_combout ),
	.datad(!\Selector3~12_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[5]~1 .extended_lut = "off";
defparam \master_writedata[5]~1 .lut_mask = 64'h0400040004000400;
defparam \master_writedata[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr5~0 (
	.dataa(!\Selector3~8_combout ),
	.datab(!\Selector11~0_combout ),
	.datac(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datad(!\master_writedata[5]~1_combout ),
	.datae(!\Selector8~0_combout ),
	.dataf(!\Selector7~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr5~0 .extended_lut = "off";
defparam \WideOr5~0 .lut_mask = 64'h333BFF7FFFFFFFFF;
defparam \WideOr5~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr17~1 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\Selector13~0_combout ),
	.datad(!\state.ST_WRITE_RECONFIG_BASIC_LCH~q ),
	.datae(!\Selector2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~1 .extended_lut = "off";
defparam \WideOr17~1 .lut_mask = 64'hF0200000F0200000;
defparam \WideOr17~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!mutex_req1),
	.datab(!\Selector1~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\WideOr6~1_combout ),
	.datae(!\WideOr5~0_combout ),
	.dataf(!\WideOr17~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'h7777777777737777;
defparam \Selector29~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr7(
	.dataa(!\WideOr7~0_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr7~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr7.extended_lut = "off";
defparam WideOr7.lut_mask = 64'h4444444444444444;
defparam WideOr7.shared_arith = "off";

cyclonev_lcell_comb WideOr6(
	.dataa(!\WideOr6~1_combout ),
	.datab(!\Selector14~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr6~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr6.extended_lut = "off";
defparam WideOr6.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam WideOr6.shared_arith = "off";

cyclonev_lcell_comb WideOr9(
	.dataa(!\Selector3~7_combout ),
	.datab(!\Selector11~0_combout ),
	.datac(!\Selector6~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr9~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr9.extended_lut = "off";
defparam WideOr9.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam WideOr9.shared_arith = "off";

cyclonev_lcell_comb \ph_readdata[13]~0 (
	.dataa(!basic_reconfig_waitrequest2),
	.datab(!\state.ST_CHECK_PHY_ADD_LEGAL~q ),
	.datac(!\state.ST_CHECK_CTRLLOCK~q ),
	.datad(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datae(!\Selector12~0_combout ),
	.dataf(!\phy_addr_is_set~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ph_readdata[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ph_readdata[13]~0 .extended_lut = "off";
defparam \ph_readdata[13]~0 .lut_mask = 64'h8C8C0088048C0088;
defparam \ph_readdata[13]~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!lif_waitrequest),
	.datab(!basic_reconfig_waitrequest1),
	.datac(!\state.ST_RELEASE_REQ~q ),
	.datad(!\Selector1~0_combout ),
	.datae(!ctrl_lock),
	.dataf(!\state.ST_CHECK_CTRLLOCK~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'hF200F2000000F200;
defparam \Selector16~0 .shared_arith = "off";

cyclonev_lcell_comb \ph_readdata[13]~1 (
	.dataa(!\Selector0~0_combout ),
	.datab(!\WideOr6~1_combout ),
	.datac(!\WideOr5~0_combout ),
	.datad(!\WideOr17~1_combout ),
	.datae(!\ph_readdata[13]~0_combout ),
	.dataf(!\Selector16~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ph_readdata[13]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ph_readdata[13]~1 .extended_lut = "off";
defparam \ph_readdata[13]~1 .lut_mask = 64'h0000000000100000;
defparam \ph_readdata[13]~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!ctrl_opcode_2),
	.datab(!ctrl_opcode_0),
	.datac(!\Selector10~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h0404040404040404;
defparam \Selector27~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~1 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(!logical_ch_addr[1]),
	.datad(!\Selector27~0_combout ),
	.datae(!ctrl_addr_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~1 .extended_lut = "off";
defparam \Selector27~1 .lut_mask = 64'hFA00C800FA00C800;
defparam \Selector27~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~2 (
	.dataa(!\Selector15~2_combout ),
	.datab(!\Selector5~2_combout ),
	.datac(!\Selector8~1_combout ),
	.datad(!ctrl_wdata_1),
	.datae(!\Selector27~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~2 .extended_lut = "off";
defparam \Selector27~2 .lut_mask = 64'hFFFF777FFFFF777F;
defparam \Selector27~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector14~0_combout ),
	.datac(!logical_ch_addr[2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \Selector26~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~1 (
	.dataa(!\Selector8~1_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(!ctrl_wdata_2),
	.datad(!ctrl_addr_5),
	.datae(!\Selector26~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~1 .extended_lut = "off";
defparam \Selector26~1 .lut_mask = 64'hFFFF0537FFFF0537;
defparam \Selector26~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector7~1_combout ),
	.datac(!logical_ch_addr[0]),
	.datad(!ctrl_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h0537053705370537;
defparam \Selector28~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~1 (
	.dataa(!\Selector5~2_combout ),
	.datab(!\Selector10~0_combout ),
	.datac(!\Selector8~1_combout ),
	.datad(!ctrl_wdata_0),
	.datae(!\Selector28~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~1 .extended_lut = "off";
defparam \Selector28~1 .lut_mask = 64'h777FFFFF777FFFFF;
defparam \Selector28~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector8~1_combout ),
	.datac(!logical_ch_addr[3]),
	.datad(!ctrl_wdata_3),
	.datae(!\Selector27~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h0537FFFF0537FFFF;
defparam \Selector25~0 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[5]~2 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector8~1_combout ),
	.datac(!\Selector7~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[5]~2 .extended_lut = "off";
defparam \master_writedata[5]~2 .lut_mask = 64'h8C8C8C8C8C8C8C8C;
defparam \master_writedata[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata[5]~3 (
	.dataa(!\Selector3~8_combout ),
	.datab(!\state.ST_WRITE_DATA_TO_RECONFIG_BASIC~q ),
	.datac(!\master_writedata[5]~1_combout ),
	.datad(!\Selector8~0_combout ),
	.datae(!\Selector7~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata[5]~3 .extended_lut = "off";
defparam \master_writedata[5]~3 .lut_mask = 64'hFD5D0000FD5D0000;
defparam \master_writedata[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!logical_ch_addr[4]),
	.datab(!ctrl_addr_4),
	.datac(!\master_writedata[5]~2_combout ),
	.datad(!\master_writedata[5]~3_combout ),
	.datae(!ctrl_wdata_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h0350F3500350F350;
defparam \Selector24~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector23~0 (
	.dataa(!logical_ch_addr[5]),
	.datab(!ctrl_addr_5),
	.datac(!\master_writedata[5]~2_combout ),
	.datad(!\master_writedata[5]~3_combout ),
	.datae(!ctrl_wdata_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h0350F3500350F350;
defparam \Selector23~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector22~0 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector8~1_combout ),
	.datac(!logical_ch_addr[6]),
	.datad(!ctrl_wdata_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector22~0 .extended_lut = "off";
defparam \Selector22~0 .lut_mask = 64'h0537053705370537;
defparam \Selector22~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector21~0 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector8~1_combout ),
	.datac(!logical_ch_addr[7]),
	.datad(!ctrl_wdata_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~0 .extended_lut = "off";
defparam \Selector21~0 .lut_mask = 64'h0537053705370537;
defparam \Selector21~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector8~1_combout ),
	.datac(!logical_ch_addr[8]),
	.datad(!ctrl_wdata_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h0537053705370537;
defparam \Selector20~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\Selector8~1_combout ),
	.datac(!logical_ch_addr[9]),
	.datad(!ctrl_wdata_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h0537053705370537;
defparam \Selector19~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h1111111111111111;
defparam \Selector18~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'h1111111111111111;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~4 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~4 .extended_lut = "off";
defparam \master_writedata~4 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~4 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~5 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~5 .extended_lut = "off";
defparam \master_writedata~5 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~5 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~6 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~6 .extended_lut = "off";
defparam \master_writedata~6 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~6 .shared_arith = "off";

cyclonev_lcell_comb \master_writedata~7 (
	.dataa(!\Selector8~1_combout ),
	.datab(!ctrl_wdata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_writedata~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_writedata~7 .extended_lut = "off";
defparam \master_writedata~7 .lut_mask = 64'h1111111111111111;
defparam \master_writedata~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~1 (
	.dataa(!\WideOr6~1_combout ),
	.datab(!\WideOr5~0_combout ),
	.datac(!\WideOr17~1_combout ),
	.datad(!\Selector16~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~1 .extended_lut = "off";
defparam \Selector16~1 .lut_mask = 64'h0004000400040004;
defparam \Selector16~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~2 (
	.dataa(!ctrl_lock),
	.datab(!\Selector4~0_combout ),
	.datac(!\Selector12~1_combout ),
	.datad(!\Selector16~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~2 .extended_lut = "off";
defparam \Selector16~2 .lut_mask = 64'hFF3BFF3BFF3BFF3B;
defparam \Selector16~2 .shared_arith = "off";

cyclonev_lcell_comb \readdata_for_user[0]~0 (
	.dataa(!\state.ST_CLR_RECONFIG_BASIC_PADDR_MODE~q ),
	.datab(!\state.ST_READ_RECONFIG_BASIC_DATA~q ),
	.datac(!\Selector12~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata_for_user[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata_for_user[0]~0 .extended_lut = "off";
defparam \readdata_for_user[0]~0 .lut_mask = 64'h0707070707070707;
defparam \readdata_for_user[0]~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xreconf_uif_2 (
	user_reconfig_readdata_10,
	user_reconfig_readdata_11,
	user_reconfig_readdata_12,
	user_reconfig_readdata_13,
	user_reconfig_readdata_14,
	user_reconfig_readdata_15,
	user_reconfig_readdata_16,
	user_reconfig_readdata_17,
	user_reconfig_readdata_18,
	user_reconfig_readdata_19,
	user_reconfig_readdata_20,
	user_reconfig_readdata_21,
	user_reconfig_readdata_22,
	user_reconfig_readdata_23,
	user_reconfig_readdata_24,
	uif_rdata_3,
	uif_rdata_4,
	uif_rdata_5,
	uif_rdata_6,
	uif_rdata_7,
	uif_rdata_8,
	uif_rdata_9,
	uif_rdata_10,
	uif_rdata_11,
	uif_rdata_12,
	uif_rdata_13,
	uif_rdata_14,
	uif_rdata_15,
	uif_rdata_16,
	uif_rdata_17,
	uif_rdata_18,
	uif_rdata_19,
	user_reconfig_readdata_0,
	Equal4,
	user_reconfig_readdata_1,
	user_reconfig_readdata_2,
	user_reconfig_readdata_3,
	user_reconfig_readdata_4,
	user_reconfig_readdata_5,
	user_reconfig_readdata_6,
	user_reconfig_readdata_7,
	user_reconfig_readdata_8,
	user_reconfig_readdata_9,
	user_reconfig_readdata_25,
	user_reconfig_readdata_26,
	user_reconfig_readdata_27,
	user_reconfig_readdata_28,
	user_reconfig_readdata_29,
	user_reconfig_readdata_30,
	user_reconfig_readdata_31,
	resync_chains0sync_r_1,
	launch_reg,
	wait_reg,
	pll_mif_busy,
	ifsel_notdone_resync,
	uif_writedata_0,
	uif_mode_1,
	uif_mode_0,
	Equal41,
	uif_rdata_0,
	ph_readdata_0,
	uif_logical_ch_addr_0,
	uif_addr_offset_0,
	comb,
	uif_writedata_1,
	uif_rdata_1,
	ph_readdata_1,
	uif_logical_ch_addr_1,
	uif_addr_offset_1,
	uif_writedata_2,
	uif_rdata_2,
	ph_readdata_2,
	uif_logical_ch_addr_2,
	uif_addr_offset_2,
	ph_readdata_3,
	uif_logical_ch_addr_3,
	user_reconfig_readdata_101,
	ph_readdata_4,
	uif_logical_ch_addr_4,
	ph_readdata_5,
	uif_logical_ch_addr_5,
	ph_readdata_6,
	uif_logical_ch_addr_6,
	ph_readdata_7,
	uif_logical_ch_addr_7,
	uif_logical_ch_addr_8,
	ph_readdata_8,
	ph_readdata_9,
	uif_logical_ch_addr_9,
	uif_addr_err,
	illegal_phy_ch,
	ph_readdata_10,
	ph_readdata_11,
	ph_readdata_12,
	ph_readdata_13,
	ph_readdata_14,
	ph_readdata_15,
	ph_readdata_16,
	ph_readdata_17,
	ph_readdata_18,
	ph_readdata_19,
	ph_readdata_20,
	uif_rdata_20,
	ph_readdata_21,
	uif_rdata_21,
	ph_readdata_22,
	uif_rdata_22,
	ph_readdata_23,
	uif_rdata_23,
	ph_readdata_24,
	uif_rdata_24,
	ph_readdata_25,
	ph_readdata_26,
	ph_readdata_27,
	ph_readdata_28,
	ph_readdata_29,
	ph_readdata_30,
	ph_readdata_31,
	uif_go1,
	uif_mode_01,
	Mux0,
	Mux3,
	WideOr0,
	reconfig_mgmt_address_1,
	reconfig_mgmt_address_0,
	reconfig_mgmt_address_2,
	reconfig_mgmt_write,
	reconfig_mgmt_read,
	mgmt_clk_clk,
	reconfig_mgmt_writedata_0,
	reconfig_mgmt_writedata_1,
	reconfig_mgmt_writedata_2,
	reconfig_mgmt_writedata_3,
	reconfig_mgmt_writedata_16,
	reconfig_mgmt_writedata_17,
	reconfig_mgmt_writedata_18,
	reconfig_mgmt_writedata_19,
	reconfig_mgmt_writedata_20,
	reconfig_mgmt_writedata_4,
	reconfig_mgmt_writedata_21,
	reconfig_mgmt_writedata_5,
	reconfig_mgmt_writedata_22,
	reconfig_mgmt_writedata_6,
	reconfig_mgmt_writedata_23,
	reconfig_mgmt_writedata_7,
	reconfig_mgmt_writedata_24,
	reconfig_mgmt_writedata_8,
	reconfig_mgmt_writedata_25,
	reconfig_mgmt_writedata_9,
	reconfig_mgmt_writedata_26,
	reconfig_mgmt_writedata_10,
	reconfig_mgmt_writedata_27,
	reconfig_mgmt_writedata_11,
	reconfig_mgmt_writedata_28,
	reconfig_mgmt_writedata_12,
	reconfig_mgmt_writedata_29,
	reconfig_mgmt_writedata_13,
	reconfig_mgmt_writedata_30,
	reconfig_mgmt_writedata_14,
	reconfig_mgmt_writedata_31,
	reconfig_mgmt_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	user_reconfig_readdata_10;
output 	user_reconfig_readdata_11;
output 	user_reconfig_readdata_12;
output 	user_reconfig_readdata_13;
output 	user_reconfig_readdata_14;
output 	user_reconfig_readdata_15;
output 	user_reconfig_readdata_16;
output 	user_reconfig_readdata_17;
output 	user_reconfig_readdata_18;
output 	user_reconfig_readdata_19;
output 	user_reconfig_readdata_20;
output 	user_reconfig_readdata_21;
output 	user_reconfig_readdata_22;
output 	user_reconfig_readdata_23;
output 	user_reconfig_readdata_24;
input 	uif_rdata_3;
input 	uif_rdata_4;
input 	uif_rdata_5;
input 	uif_rdata_6;
input 	uif_rdata_7;
input 	uif_rdata_8;
input 	uif_rdata_9;
input 	uif_rdata_10;
input 	uif_rdata_11;
input 	uif_rdata_12;
input 	uif_rdata_13;
input 	uif_rdata_14;
input 	uif_rdata_15;
input 	uif_rdata_16;
input 	uif_rdata_17;
input 	uif_rdata_18;
input 	uif_rdata_19;
output 	user_reconfig_readdata_0;
input 	Equal4;
output 	user_reconfig_readdata_1;
output 	user_reconfig_readdata_2;
output 	user_reconfig_readdata_3;
output 	user_reconfig_readdata_4;
output 	user_reconfig_readdata_5;
output 	user_reconfig_readdata_6;
output 	user_reconfig_readdata_7;
output 	user_reconfig_readdata_8;
output 	user_reconfig_readdata_9;
output 	user_reconfig_readdata_25;
output 	user_reconfig_readdata_26;
output 	user_reconfig_readdata_27;
output 	user_reconfig_readdata_28;
output 	user_reconfig_readdata_29;
output 	user_reconfig_readdata_30;
output 	user_reconfig_readdata_31;
output 	resync_chains0sync_r_1;
output 	launch_reg;
output 	wait_reg;
input 	pll_mif_busy;
input 	ifsel_notdone_resync;
output 	uif_writedata_0;
output 	uif_mode_1;
output 	uif_mode_0;
input 	Equal41;
input 	uif_rdata_0;
input 	ph_readdata_0;
output 	uif_logical_ch_addr_0;
output 	uif_addr_offset_0;
input 	comb;
output 	uif_writedata_1;
input 	uif_rdata_1;
input 	ph_readdata_1;
output 	uif_logical_ch_addr_1;
output 	uif_addr_offset_1;
output 	uif_writedata_2;
input 	uif_rdata_2;
input 	ph_readdata_2;
output 	uif_logical_ch_addr_2;
output 	uif_addr_offset_2;
input 	ph_readdata_3;
output 	uif_logical_ch_addr_3;
output 	user_reconfig_readdata_101;
input 	ph_readdata_4;
output 	uif_logical_ch_addr_4;
input 	ph_readdata_5;
output 	uif_logical_ch_addr_5;
input 	ph_readdata_6;
output 	uif_logical_ch_addr_6;
input 	ph_readdata_7;
output 	uif_logical_ch_addr_7;
output 	uif_logical_ch_addr_8;
input 	ph_readdata_8;
input 	ph_readdata_9;
output 	uif_logical_ch_addr_9;
input 	uif_addr_err;
input 	illegal_phy_ch;
input 	ph_readdata_10;
input 	ph_readdata_11;
input 	ph_readdata_12;
input 	ph_readdata_13;
input 	ph_readdata_14;
input 	ph_readdata_15;
input 	ph_readdata_16;
input 	ph_readdata_17;
input 	ph_readdata_18;
input 	ph_readdata_19;
input 	ph_readdata_20;
input 	uif_rdata_20;
input 	ph_readdata_21;
input 	uif_rdata_21;
input 	ph_readdata_22;
input 	uif_rdata_22;
input 	ph_readdata_23;
input 	uif_rdata_23;
input 	ph_readdata_24;
input 	uif_rdata_24;
input 	ph_readdata_25;
input 	ph_readdata_26;
input 	ph_readdata_27;
input 	ph_readdata_28;
input 	ph_readdata_29;
input 	ph_readdata_30;
input 	ph_readdata_31;
output 	uif_go1;
input 	uif_mode_01;
output 	Mux0;
output 	Mux3;
input 	WideOr0;
input 	reconfig_mgmt_address_1;
input 	reconfig_mgmt_address_0;
input 	reconfig_mgmt_address_2;
input 	reconfig_mgmt_write;
input 	reconfig_mgmt_read;
input 	mgmt_clk_clk;
input 	reconfig_mgmt_writedata_0;
input 	reconfig_mgmt_writedata_1;
input 	reconfig_mgmt_writedata_2;
input 	reconfig_mgmt_writedata_3;
input 	reconfig_mgmt_writedata_16;
input 	reconfig_mgmt_writedata_17;
input 	reconfig_mgmt_writedata_18;
input 	reconfig_mgmt_writedata_19;
input 	reconfig_mgmt_writedata_20;
input 	reconfig_mgmt_writedata_4;
input 	reconfig_mgmt_writedata_21;
input 	reconfig_mgmt_writedata_5;
input 	reconfig_mgmt_writedata_22;
input 	reconfig_mgmt_writedata_6;
input 	reconfig_mgmt_writedata_23;
input 	reconfig_mgmt_writedata_7;
input 	reconfig_mgmt_writedata_24;
input 	reconfig_mgmt_writedata_8;
input 	reconfig_mgmt_writedata_25;
input 	reconfig_mgmt_writedata_9;
input 	reconfig_mgmt_writedata_26;
input 	reconfig_mgmt_writedata_10;
input 	reconfig_mgmt_writedata_27;
input 	reconfig_mgmt_writedata_11;
input 	reconfig_mgmt_writedata_28;
input 	reconfig_mgmt_writedata_12;
input 	reconfig_mgmt_writedata_29;
input 	reconfig_mgmt_writedata_13;
input 	reconfig_mgmt_writedata_30;
input 	reconfig_mgmt_writedata_14;
input 	reconfig_mgmt_writedata_31;
input 	reconfig_mgmt_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \uif_writedata[0]~0_combout ;
wire \uif_writedata[10]~q ;
wire \Mux25~0_combout ;
wire \user_reconfig_readdata[3]~8_combout ;
wire \uif_writedata[11]~q ;
wire \Mux24~0_combout ;
wire \uif_writedata[12]~q ;
wire \Mux23~0_combout ;
wire \uif_writedata[13]~q ;
wire \Mux22~0_combout ;
wire \uif_writedata[14]~q ;
wire \Mux21~0_combout ;
wire \uif_writedata[15]~q ;
wire \Mux20~0_combout ;
wire \uif_writedata[16]~q ;
wire \Mux19~0_combout ;
wire \uif_writedata[17]~q ;
wire \Mux18~0_combout ;
wire \uif_writedata[18]~q ;
wire \Mux17~0_combout ;
wire \uif_writedata[19]~q ;
wire \Mux16~0_combout ;
wire \uif_writedata[20]~q ;
wire \Mux15~0_combout ;
wire \uif_writedata[21]~q ;
wire \Mux14~0_combout ;
wire \uif_writedata[22]~q ;
wire \Mux13~0_combout ;
wire \uif_writedata[23]~q ;
wire \Mux12~0_combout ;
wire \uif_writedata[24]~q ;
wire \Mux11~0_combout ;
wire \user_reconfig_readdata[2]~0_combout ;
wire \user_reconfig_readdata[2]~1_combout ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \user_reconfig_readdata[0]~2_combout ;
wire \user_reconfig_readdata[0]~3_combout ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \user_reconfig_readdata[3]~4_combout ;
wire \Mux32~0_combout ;
wire \user_reconfig_readdata[3]~5_combout ;
wire \user_reconfig_readdata[3]~6_combout ;
wire \uif_writedata[3]~q ;
wire \Mux32~1_combout ;
wire \Mux32~2_combout ;
wire \uif_writedata[4]~q ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \uif_writedata[5]~q ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \uif_writedata[6]~q ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \uif_writedata[7]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \uif_writedata[8]~q ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \uif_writedata[9]~q ;
wire \illegal_addr_error~0_combout ;
wire \illegal_addr_error~q ;
wire \Mux26~1_combout ;
wire \Mux26~0_combout ;
wire \user_reconfig_readdata[27]~9_combout ;
wire \uif_writedata[25]~q ;
wire \Mux10~0_combout ;
wire \uif_writedata[26]~q ;
wire \Mux9~0_combout ;
wire \uif_writedata[27]~q ;
wire \Mux8~0_combout ;
wire \uif_writedata[28]~q ;
wire \Mux7~0_combout ;
wire \uif_writedata[29]~q ;
wire \Mux6~0_combout ;
wire \uif_writedata[30]~q ;
wire \Mux5~0_combout ;
wire \uif_writedata[31]~q ;
wire \Mux4~0_combout ;
wire \uif_mode[1]~1_combout ;
wire \Mux0~1_combout ;
wire \uif_mode[0]~0_combout ;
wire \uif_logical_ch_addr[0]~0_combout ;
wire \uif_addr_offset[2]~0_combout ;
wire \Mux0~2_combout ;


RECONFIGURE_IP_altera_wait_generate_3 wait_gen(
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.launch_reg1(launch_reg),
	.wait_reg1(wait_reg),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.launch_signal(comb),
	.mgmt_clk_clk(mgmt_clk_clk));

dffeas \user_reconfig_readdata[10] (
	.clk(mgmt_clk_clk),
	.d(\Mux25~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_10),
	.prn(vcc));
defparam \user_reconfig_readdata[10] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[10] .power_up = "low";

dffeas \user_reconfig_readdata[11] (
	.clk(mgmt_clk_clk),
	.d(\Mux24~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_11),
	.prn(vcc));
defparam \user_reconfig_readdata[11] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[11] .power_up = "low";

dffeas \user_reconfig_readdata[12] (
	.clk(mgmt_clk_clk),
	.d(\Mux23~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_12),
	.prn(vcc));
defparam \user_reconfig_readdata[12] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[12] .power_up = "low";

dffeas \user_reconfig_readdata[13] (
	.clk(mgmt_clk_clk),
	.d(\Mux22~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_13),
	.prn(vcc));
defparam \user_reconfig_readdata[13] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[13] .power_up = "low";

dffeas \user_reconfig_readdata[14] (
	.clk(mgmt_clk_clk),
	.d(\Mux21~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_14),
	.prn(vcc));
defparam \user_reconfig_readdata[14] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[14] .power_up = "low";

dffeas \user_reconfig_readdata[15] (
	.clk(mgmt_clk_clk),
	.d(\Mux20~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_15),
	.prn(vcc));
defparam \user_reconfig_readdata[15] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[15] .power_up = "low";

dffeas \user_reconfig_readdata[16] (
	.clk(mgmt_clk_clk),
	.d(\Mux19~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_16),
	.prn(vcc));
defparam \user_reconfig_readdata[16] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[16] .power_up = "low";

dffeas \user_reconfig_readdata[17] (
	.clk(mgmt_clk_clk),
	.d(\Mux18~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_17),
	.prn(vcc));
defparam \user_reconfig_readdata[17] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[17] .power_up = "low";

dffeas \user_reconfig_readdata[18] (
	.clk(mgmt_clk_clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_18),
	.prn(vcc));
defparam \user_reconfig_readdata[18] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[18] .power_up = "low";

dffeas \user_reconfig_readdata[19] (
	.clk(mgmt_clk_clk),
	.d(\Mux16~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_19),
	.prn(vcc));
defparam \user_reconfig_readdata[19] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[19] .power_up = "low";

dffeas \user_reconfig_readdata[20] (
	.clk(mgmt_clk_clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_20),
	.prn(vcc));
defparam \user_reconfig_readdata[20] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[20] .power_up = "low";

dffeas \user_reconfig_readdata[21] (
	.clk(mgmt_clk_clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_21),
	.prn(vcc));
defparam \user_reconfig_readdata[21] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[21] .power_up = "low";

dffeas \user_reconfig_readdata[22] (
	.clk(mgmt_clk_clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_22),
	.prn(vcc));
defparam \user_reconfig_readdata[22] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[22] .power_up = "low";

dffeas \user_reconfig_readdata[23] (
	.clk(mgmt_clk_clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_23),
	.prn(vcc));
defparam \user_reconfig_readdata[23] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[23] .power_up = "low";

dffeas \user_reconfig_readdata[24] (
	.clk(mgmt_clk_clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(user_reconfig_readdata_101),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_24),
	.prn(vcc));
defparam \user_reconfig_readdata[24] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[24] .power_up = "low";

dffeas \user_reconfig_readdata[0] (
	.clk(mgmt_clk_clk),
	.d(\Mux35~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_0),
	.prn(vcc));
defparam \user_reconfig_readdata[0] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[0] .power_up = "low";

dffeas \user_reconfig_readdata[1] (
	.clk(mgmt_clk_clk),
	.d(\Mux34~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_1),
	.prn(vcc));
defparam \user_reconfig_readdata[1] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[1] .power_up = "low";

dffeas \user_reconfig_readdata[2] (
	.clk(mgmt_clk_clk),
	.d(\Mux33~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_2),
	.prn(vcc));
defparam \user_reconfig_readdata[2] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[2] .power_up = "low";

dffeas \user_reconfig_readdata[3] (
	.clk(mgmt_clk_clk),
	.d(\Mux32~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_3),
	.prn(vcc));
defparam \user_reconfig_readdata[3] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[3] .power_up = "low";

dffeas \user_reconfig_readdata[4] (
	.clk(mgmt_clk_clk),
	.d(\Mux31~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_4),
	.prn(vcc));
defparam \user_reconfig_readdata[4] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[4] .power_up = "low";

dffeas \user_reconfig_readdata[5] (
	.clk(mgmt_clk_clk),
	.d(\Mux30~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_5),
	.prn(vcc));
defparam \user_reconfig_readdata[5] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[5] .power_up = "low";

dffeas \user_reconfig_readdata[6] (
	.clk(mgmt_clk_clk),
	.d(\Mux29~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_6),
	.prn(vcc));
defparam \user_reconfig_readdata[6] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[6] .power_up = "low";

dffeas \user_reconfig_readdata[7] (
	.clk(mgmt_clk_clk),
	.d(\Mux28~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_7),
	.prn(vcc));
defparam \user_reconfig_readdata[7] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[7] .power_up = "low";

dffeas \user_reconfig_readdata[8] (
	.clk(mgmt_clk_clk),
	.d(\Mux27~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_8),
	.prn(vcc));
defparam \user_reconfig_readdata[8] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[8] .power_up = "low";

dffeas \user_reconfig_readdata[9] (
	.clk(mgmt_clk_clk),
	.d(\Mux26~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[0]~3_combout ),
	.q(user_reconfig_readdata_9),
	.prn(vcc));
defparam \user_reconfig_readdata[9] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[9] .power_up = "low";

dffeas \user_reconfig_readdata[25] (
	.clk(mgmt_clk_clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_25),
	.prn(vcc));
defparam \user_reconfig_readdata[25] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[25] .power_up = "low";

dffeas \user_reconfig_readdata[26] (
	.clk(mgmt_clk_clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_26),
	.prn(vcc));
defparam \user_reconfig_readdata[26] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[26] .power_up = "low";

dffeas \user_reconfig_readdata[27] (
	.clk(mgmt_clk_clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_27),
	.prn(vcc));
defparam \user_reconfig_readdata[27] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[27] .power_up = "low";

dffeas \user_reconfig_readdata[28] (
	.clk(mgmt_clk_clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_28),
	.prn(vcc));
defparam \user_reconfig_readdata[28] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[28] .power_up = "low";

dffeas \user_reconfig_readdata[29] (
	.clk(mgmt_clk_clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_29),
	.prn(vcc));
defparam \user_reconfig_readdata[29] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[29] .power_up = "low";

dffeas \user_reconfig_readdata[30] (
	.clk(mgmt_clk_clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_30),
	.prn(vcc));
defparam \user_reconfig_readdata[30] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[30] .power_up = "low";

dffeas \user_reconfig_readdata[31] (
	.clk(mgmt_clk_clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\user_reconfig_readdata[3]~8_combout ),
	.q(user_reconfig_readdata_31),
	.prn(vcc));
defparam \user_reconfig_readdata[31] .is_wysiwyg = "true";
defparam \user_reconfig_readdata[31] .power_up = "low";

dffeas \uif_writedata[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_0),
	.prn(vcc));
defparam \uif_writedata[0] .is_wysiwyg = "true";
defparam \uif_writedata[0] .power_up = "low";

dffeas \uif_mode[1] (
	.clk(mgmt_clk_clk),
	.d(\uif_mode[1]~1_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_mode[0]~0_combout ),
	.q(uif_mode_1),
	.prn(vcc));
defparam \uif_mode[1] .is_wysiwyg = "true";
defparam \uif_mode[1] .power_up = "low";

dffeas \uif_mode[0] (
	.clk(mgmt_clk_clk),
	.d(Mux3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_mode[0]~0_combout ),
	.q(uif_mode_0),
	.prn(vcc));
defparam \uif_mode[0] .is_wysiwyg = "true";
defparam \uif_mode[0] .power_up = "low";

dffeas \uif_logical_ch_addr[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_0),
	.prn(vcc));
defparam \uif_logical_ch_addr[0] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[0] .power_up = "low";

dffeas \uif_addr_offset[0] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_0),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[2]~0_combout ),
	.q(uif_addr_offset_0),
	.prn(vcc));
defparam \uif_addr_offset[0] .is_wysiwyg = "true";
defparam \uif_addr_offset[0] .power_up = "low";

dffeas \uif_writedata[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_1),
	.prn(vcc));
defparam \uif_writedata[1] .is_wysiwyg = "true";
defparam \uif_writedata[1] .power_up = "low";

dffeas \uif_logical_ch_addr[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_1),
	.prn(vcc));
defparam \uif_logical_ch_addr[1] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[1] .power_up = "low";

dffeas \uif_addr_offset[1] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_1),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[2]~0_combout ),
	.q(uif_addr_offset_1),
	.prn(vcc));
defparam \uif_addr_offset[1] .is_wysiwyg = "true";
defparam \uif_addr_offset[1] .power_up = "low";

dffeas \uif_writedata[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(uif_writedata_2),
	.prn(vcc));
defparam \uif_writedata[2] .is_wysiwyg = "true";
defparam \uif_writedata[2] .power_up = "low";

dffeas \uif_logical_ch_addr[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_2),
	.prn(vcc));
defparam \uif_logical_ch_addr[2] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[2] .power_up = "low";

dffeas \uif_addr_offset[2] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_2),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_addr_offset[2]~0_combout ),
	.q(uif_addr_offset_2),
	.prn(vcc));
defparam \uif_addr_offset[2] .is_wysiwyg = "true";
defparam \uif_addr_offset[2] .power_up = "low";

dffeas \uif_logical_ch_addr[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_3),
	.prn(vcc));
defparam \uif_logical_ch_addr[3] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[3] .power_up = "low";

cyclonev_lcell_comb \user_reconfig_readdata[10]~7 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(user_reconfig_readdata_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[10]~7 .extended_lut = "off";
defparam \user_reconfig_readdata[10]~7 .lut_mask = 64'hD7D7D7D7D7D7D7D7;
defparam \user_reconfig_readdata[10]~7 .shared_arith = "off";

dffeas \uif_logical_ch_addr[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_4),
	.prn(vcc));
defparam \uif_logical_ch_addr[4] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[4] .power_up = "low";

dffeas \uif_logical_ch_addr[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_5),
	.prn(vcc));
defparam \uif_logical_ch_addr[5] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[5] .power_up = "low";

dffeas \uif_logical_ch_addr[6] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_6),
	.prn(vcc));
defparam \uif_logical_ch_addr[6] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[6] .power_up = "low";

dffeas \uif_logical_ch_addr[7] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_7),
	.prn(vcc));
defparam \uif_logical_ch_addr[7] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[7] .power_up = "low";

dffeas \uif_logical_ch_addr[8] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_8),
	.prn(vcc));
defparam \uif_logical_ch_addr[8] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[8] .power_up = "low";

dffeas \uif_logical_ch_addr[9] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_logical_ch_addr[0]~0_combout ),
	.q(uif_logical_ch_addr_9),
	.prn(vcc));
defparam \uif_logical_ch_addr[9] .is_wysiwyg = "true";
defparam \uif_logical_ch_addr[9] .power_up = "low";

dffeas uif_go(
	.clk(mgmt_clk_clk),
	.d(\Mux0~2_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_go1),
	.prn(vcc));
defparam uif_go.is_wysiwyg = "true";
defparam uif_go.power_up = "low";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h6060606060606060;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_writedata_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h1111111111111111;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!Equal4),
	.datab(!reconfig_mgmt_write),
	.datac(!pll_mif_busy),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h1010101010101010;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_writedata[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_writedata[0]~0 .extended_lut = "off";
defparam \uif_writedata[0]~0 .lut_mask = 64'h0008000800080008;
defparam \uif_writedata[0]~0 .shared_arith = "off";

dffeas \uif_writedata[10] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_10),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[10]~q ),
	.prn(vcc));
defparam \uif_writedata[10] .is_wysiwyg = "true";
defparam \uif_writedata[10] .power_up = "low";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_10),
	.datad(!\uif_writedata[10]~q ),
	.datae(!uif_rdata_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "off";
defparam \Mux25~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[3]~8 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!comb),
	.datac(!pll_mif_busy),
	.datad(!uif_mode_1),
	.datae(!uif_mode_0),
	.dataf(!user_reconfig_readdata_101),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[3]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[3]~8 .extended_lut = "off";
defparam \user_reconfig_readdata[3]~8 .lut_mask = 64'h3030302033333333;
defparam \user_reconfig_readdata[3]~8 .shared_arith = "off";

dffeas \uif_writedata[11] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_11),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[11]~q ),
	.prn(vcc));
defparam \uif_writedata[11] .is_wysiwyg = "true";
defparam \uif_writedata[11] .power_up = "low";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_11),
	.datad(!\uif_writedata[11]~q ),
	.datae(!uif_rdata_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "off";
defparam \Mux24~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux24~0 .shared_arith = "off";

dffeas \uif_writedata[12] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_12),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[12]~q ),
	.prn(vcc));
defparam \uif_writedata[12] .is_wysiwyg = "true";
defparam \uif_writedata[12] .power_up = "low";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_12),
	.datad(!\uif_writedata[12]~q ),
	.datae(!uif_rdata_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "off";
defparam \Mux23~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux23~0 .shared_arith = "off";

dffeas \uif_writedata[13] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_13),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[13]~q ),
	.prn(vcc));
defparam \uif_writedata[13] .is_wysiwyg = "true";
defparam \uif_writedata[13] .power_up = "low";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_13),
	.datad(!\uif_writedata[13]~q ),
	.datae(!uif_rdata_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "off";
defparam \Mux22~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux22~0 .shared_arith = "off";

dffeas \uif_writedata[14] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_14),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[14]~q ),
	.prn(vcc));
defparam \uif_writedata[14] .is_wysiwyg = "true";
defparam \uif_writedata[14] .power_up = "low";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_14),
	.datad(!\uif_writedata[14]~q ),
	.datae(!uif_rdata_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "off";
defparam \Mux21~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux21~0 .shared_arith = "off";

dffeas \uif_writedata[15] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_15),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[15]~q ),
	.prn(vcc));
defparam \uif_writedata[15] .is_wysiwyg = "true";
defparam \uif_writedata[15] .power_up = "low";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_15),
	.datad(!\uif_writedata[15]~q ),
	.datae(!uif_rdata_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "off";
defparam \Mux20~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux20~0 .shared_arith = "off";

dffeas \uif_writedata[16] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_16),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[16]~q ),
	.prn(vcc));
defparam \uif_writedata[16] .is_wysiwyg = "true";
defparam \uif_writedata[16] .power_up = "low";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_16),
	.datad(!\uif_writedata[16]~q ),
	.datae(!uif_rdata_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "off";
defparam \Mux19~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux19~0 .shared_arith = "off";

dffeas \uif_writedata[17] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_17),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[17]~q ),
	.prn(vcc));
defparam \uif_writedata[17] .is_wysiwyg = "true";
defparam \uif_writedata[17] .power_up = "low";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_17),
	.datad(!\uif_writedata[17]~q ),
	.datae(!uif_rdata_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "off";
defparam \Mux18~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux18~0 .shared_arith = "off";

dffeas \uif_writedata[18] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_18),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[18]~q ),
	.prn(vcc));
defparam \uif_writedata[18] .is_wysiwyg = "true";
defparam \uif_writedata[18] .power_up = "low";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_18),
	.datad(!\uif_writedata[18]~q ),
	.datae(!uif_rdata_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "off";
defparam \Mux17~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux17~0 .shared_arith = "off";

dffeas \uif_writedata[19] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_19),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[19]~q ),
	.prn(vcc));
defparam \uif_writedata[19] .is_wysiwyg = "true";
defparam \uif_writedata[19] .power_up = "low";

cyclonev_lcell_comb \Mux16~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_19),
	.datad(!\uif_writedata[19]~q ),
	.datae(!uif_rdata_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "off";
defparam \Mux16~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux16~0 .shared_arith = "off";

dffeas \uif_writedata[20] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_20),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[20]~q ),
	.prn(vcc));
defparam \uif_writedata[20] .is_wysiwyg = "true";
defparam \uif_writedata[20] .power_up = "low";

cyclonev_lcell_comb \Mux15~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_20),
	.datad(!\uif_writedata[20]~q ),
	.datae(!uif_rdata_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~0 .extended_lut = "off";
defparam \Mux15~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux15~0 .shared_arith = "off";

dffeas \uif_writedata[21] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_21),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[21]~q ),
	.prn(vcc));
defparam \uif_writedata[21] .is_wysiwyg = "true";
defparam \uif_writedata[21] .power_up = "low";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_21),
	.datad(!\uif_writedata[21]~q ),
	.datae(!uif_rdata_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "off";
defparam \Mux14~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux14~0 .shared_arith = "off";

dffeas \uif_writedata[22] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_22),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[22]~q ),
	.prn(vcc));
defparam \uif_writedata[22] .is_wysiwyg = "true";
defparam \uif_writedata[22] .power_up = "low";

cyclonev_lcell_comb \Mux13~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_22),
	.datad(!\uif_writedata[22]~q ),
	.datae(!uif_rdata_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "off";
defparam \Mux13~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux13~0 .shared_arith = "off";

dffeas \uif_writedata[23] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_23),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[23]~q ),
	.prn(vcc));
defparam \uif_writedata[23] .is_wysiwyg = "true";
defparam \uif_writedata[23] .power_up = "low";

cyclonev_lcell_comb \Mux12~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_23),
	.datad(!\uif_writedata[23]~q ),
	.datae(!uif_rdata_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "off";
defparam \Mux12~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux12~0 .shared_arith = "off";

dffeas \uif_writedata[24] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_24),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[24]~q ),
	.prn(vcc));
defparam \uif_writedata[24] .is_wysiwyg = "true";
defparam \uif_writedata[24] .power_up = "low";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!Equal41),
	.datac(!ph_readdata_24),
	.datad(!\uif_writedata[24]~q ),
	.datae(!uif_rdata_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "off";
defparam \Mux11~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[2]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[2]~0 .extended_lut = "off";
defparam \user_reconfig_readdata[2]~0 .lut_mask = 64'h070F070F070F070F;
defparam \user_reconfig_readdata[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[2]~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[2]~1 .extended_lut = "off";
defparam \user_reconfig_readdata[2]~1 .lut_mask = 64'h0F070F070F070F07;
defparam \user_reconfig_readdata[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_0),
	.datad(!uif_logical_ch_addr_0),
	.datae(!uif_addr_offset_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~0 .extended_lut = "off";
defparam \Mux35~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux35~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~1 (
	.dataa(!uif_writedata_0),
	.datab(!\user_reconfig_readdata[2]~0_combout ),
	.datac(!\user_reconfig_readdata[2]~1_combout ),
	.datad(!uif_rdata_0),
	.datae(!\Mux35~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux35~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~1 .extended_lut = "off";
defparam \Mux35~1 .lut_mask = 64'h101CD0DC101CD0DC;
defparam \Mux35~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~2 (
	.dataa(!reconfig_mgmt_address_0),
	.datab(!pll_mif_busy),
	.datac(!uif_mode_1),
	.datad(!uif_mode_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~2 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~2 .lut_mask = 64'hCCC4CCC4CCC4CCC4;
defparam \user_reconfig_readdata[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[0]~3 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!comb),
	.datae(!\user_reconfig_readdata[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[0]~3 .extended_lut = "off";
defparam \user_reconfig_readdata[0]~3 .lut_mask = 64'h00D700FF00D700FF;
defparam \user_reconfig_readdata[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_1),
	.datad(!uif_logical_ch_addr_1),
	.datae(!uif_addr_offset_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~0 .extended_lut = "off";
defparam \Mux34~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux34~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~1 (
	.dataa(!\user_reconfig_readdata[2]~0_combout ),
	.datab(!\user_reconfig_readdata[2]~1_combout ),
	.datac(!uif_writedata_1),
	.datad(!uif_rdata_1),
	.datae(!\Mux34~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux34~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~1 .extended_lut = "off";
defparam \Mux34~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux34~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!ph_readdata_2),
	.datad(!uif_logical_ch_addr_2),
	.datae(!uif_addr_offset_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~0 .extended_lut = "off";
defparam \Mux33~0 .lut_mask = 64'h028A139B028A139B;
defparam \Mux33~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~1 (
	.dataa(!\user_reconfig_readdata[2]~0_combout ),
	.datab(!\user_reconfig_readdata[2]~1_combout ),
	.datac(!uif_writedata_2),
	.datad(!uif_rdata_2),
	.datae(!\Mux33~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux33~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~1 .extended_lut = "off";
defparam \Mux33~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux33~1 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[3]~4 (
	.dataa(!reconfig_mgmt_address_0),
	.datab(!reconfig_mgmt_address_2),
	.datac(!Equal41),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[3]~4 .extended_lut = "off";
defparam \user_reconfig_readdata[3]~4 .lut_mask = 64'h3131313131313131;
defparam \user_reconfig_readdata[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~0 .extended_lut = "off";
defparam \Mux32~0 .lut_mask = 64'h2820282028202820;
defparam \Mux32~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[3]~5 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[3]~5 .extended_lut = "off";
defparam \user_reconfig_readdata[3]~5 .lut_mask = 64'hAAA2AAA2AAA2AAA2;
defparam \user_reconfig_readdata[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[3]~6 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[3]~6 .extended_lut = "off";
defparam \user_reconfig_readdata[3]~6 .lut_mask = 64'h8088808880888088;
defparam \user_reconfig_readdata[3]~6 .shared_arith = "off";

dffeas \uif_writedata[3] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_3),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[3]~q ),
	.prn(vcc));
defparam \uif_writedata[3] .is_wysiwyg = "true";
defparam \uif_writedata[3] .power_up = "low";

cyclonev_lcell_comb \Mux32~1 (
	.dataa(!\user_reconfig_readdata[3]~5_combout ),
	.datab(!\user_reconfig_readdata[3]~6_combout ),
	.datac(!uif_logical_ch_addr_3),
	.datad(!\uif_writedata[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~1 .extended_lut = "off";
defparam \Mux32~1 .lut_mask = 64'h0123012301230123;
defparam \Mux32~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~2 (
	.dataa(!uif_rdata_3),
	.datab(!\user_reconfig_readdata[3]~4_combout ),
	.datac(!ph_readdata_3),
	.datad(!\Mux32~0_combout ),
	.datae(!\Mux32~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~2 .extended_lut = "off";
defparam \Mux32~2 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \Mux32~2 .shared_arith = "off";

dffeas \uif_writedata[4] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_4),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[4]~q ),
	.prn(vcc));
defparam \uif_writedata[4] .is_wysiwyg = "true";
defparam \uif_writedata[4] .power_up = "low";

cyclonev_lcell_comb \Mux31~0 (
	.dataa(!\user_reconfig_readdata[3]~5_combout ),
	.datab(!\user_reconfig_readdata[3]~6_combout ),
	.datac(!uif_logical_ch_addr_4),
	.datad(!\uif_writedata[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~0 .extended_lut = "off";
defparam \Mux31~0 .lut_mask = 64'h0123012301230123;
defparam \Mux31~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux31~1 (
	.dataa(!\user_reconfig_readdata[3]~4_combout ),
	.datab(!\Mux32~0_combout ),
	.datac(!uif_rdata_4),
	.datad(!ph_readdata_4),
	.datae(!\Mux31~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux31~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~1 .extended_lut = "off";
defparam \Mux31~1 .lut_mask = 64'h0123FFFF0123FFFF;
defparam \Mux31~1 .shared_arith = "off";

dffeas \uif_writedata[5] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_5),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[5]~q ),
	.prn(vcc));
defparam \uif_writedata[5] .is_wysiwyg = "true";
defparam \uif_writedata[5] .power_up = "low";

cyclonev_lcell_comb \Mux30~0 (
	.dataa(!\user_reconfig_readdata[3]~5_combout ),
	.datab(!\user_reconfig_readdata[3]~6_combout ),
	.datac(!uif_logical_ch_addr_5),
	.datad(!\uif_writedata[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~0 .extended_lut = "off";
defparam \Mux30~0 .lut_mask = 64'h0123012301230123;
defparam \Mux30~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux30~1 (
	.dataa(!\user_reconfig_readdata[3]~4_combout ),
	.datab(!\Mux32~0_combout ),
	.datac(!uif_rdata_5),
	.datad(!ph_readdata_5),
	.datae(!\Mux30~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux30~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~1 .extended_lut = "off";
defparam \Mux30~1 .lut_mask = 64'h0123FFFF0123FFFF;
defparam \Mux30~1 .shared_arith = "off";

dffeas \uif_writedata[6] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_6),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[6]~q ),
	.prn(vcc));
defparam \uif_writedata[6] .is_wysiwyg = "true";
defparam \uif_writedata[6] .power_up = "low";

cyclonev_lcell_comb \Mux29~0 (
	.dataa(!\user_reconfig_readdata[3]~5_combout ),
	.datab(!\user_reconfig_readdata[3]~6_combout ),
	.datac(!uif_logical_ch_addr_6),
	.datad(!\uif_writedata[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~0 .extended_lut = "off";
defparam \Mux29~0 .lut_mask = 64'h0123012301230123;
defparam \Mux29~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux29~1 (
	.dataa(!\user_reconfig_readdata[3]~4_combout ),
	.datab(!\Mux32~0_combout ),
	.datac(!uif_rdata_6),
	.datad(!ph_readdata_6),
	.datae(!\Mux29~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux29~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~1 .extended_lut = "off";
defparam \Mux29~1 .lut_mask = 64'h0123FFFF0123FFFF;
defparam \Mux29~1 .shared_arith = "off";

dffeas \uif_writedata[7] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_7),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[7]~q ),
	.prn(vcc));
defparam \uif_writedata[7] .is_wysiwyg = "true";
defparam \uif_writedata[7] .power_up = "low";

cyclonev_lcell_comb \Mux28~0 (
	.dataa(!\user_reconfig_readdata[3]~5_combout ),
	.datab(!\user_reconfig_readdata[3]~6_combout ),
	.datac(!uif_logical_ch_addr_7),
	.datad(!\uif_writedata[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~0 .extended_lut = "off";
defparam \Mux28~0 .lut_mask = 64'h0123012301230123;
defparam \Mux28~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~1 (
	.dataa(!\user_reconfig_readdata[3]~4_combout ),
	.datab(!\Mux32~0_combout ),
	.datac(!uif_rdata_7),
	.datad(!ph_readdata_7),
	.datae(!\Mux28~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~1 .extended_lut = "off";
defparam \Mux28~1 .lut_mask = 64'h0123FFFF0123FFFF;
defparam \Mux28~1 .shared_arith = "off";

dffeas \uif_writedata[8] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_8),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[8]~q ),
	.prn(vcc));
defparam \uif_writedata[8] .is_wysiwyg = "true";
defparam \uif_writedata[8] .power_up = "low";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!pll_mif_busy),
	.datad(!uif_logical_ch_addr_8),
	.datae(!ph_readdata_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "off";
defparam \Mux27~0 .lut_mask = 64'h048C26AE048C26AE;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~1 (
	.dataa(!\user_reconfig_readdata[2]~0_combout ),
	.datab(!\user_reconfig_readdata[2]~1_combout ),
	.datac(!\uif_writedata[8]~q ),
	.datad(!uif_rdata_8),
	.datae(!\Mux27~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~1 .extended_lut = "off";
defparam \Mux27~1 .lut_mask = 64'h04268CAE04268CAE;
defparam \Mux27~1 .shared_arith = "off";

dffeas \uif_writedata[9] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_9),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[9]~q ),
	.prn(vcc));
defparam \uif_writedata[9] .is_wysiwyg = "true";
defparam \uif_writedata[9] .power_up = "low";

cyclonev_lcell_comb \illegal_addr_error~0 (
	.dataa(!Equal4),
	.datab(!reconfig_mgmt_read),
	.datac(!reconfig_mgmt_write),
	.datad(!\illegal_addr_error~q ),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\illegal_addr_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \illegal_addr_error~0 .extended_lut = "off";
defparam \illegal_addr_error~0 .lut_mask = 64'h000015FF000015FF;
defparam \illegal_addr_error~0 .shared_arith = "off";

dffeas illegal_addr_error(
	.clk(mgmt_clk_clk),
	.d(\illegal_addr_error~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\illegal_addr_error~q ),
	.prn(vcc));
defparam illegal_addr_error.is_wysiwyg = "true";
defparam illegal_addr_error.power_up = "low";

cyclonev_lcell_comb \Mux26~1 (
	.dataa(!illegal_phy_ch),
	.datab(!uif_addr_err),
	.datac(!ph_readdata_9),
	.datad(!\illegal_addr_error~q ),
	.datae(!reconfig_mgmt_address_0),
	.dataf(!reconfig_mgmt_address_1),
	.datag(!uif_logical_ch_addr_9),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~1 .extended_lut = "on";
defparam \Mux26~1 .lut_mask = 64'h0F0F0F0F77FF0000;
defparam \Mux26~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!\user_reconfig_readdata[2]~0_combout ),
	.datab(!\user_reconfig_readdata[2]~1_combout ),
	.datac(!\uif_writedata[9]~q ),
	.datad(!\Mux26~1_combout ),
	.datae(!uif_rdata_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "off";
defparam \Mux26~0 .lut_mask = 64'h048C26AE048C26AE;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \user_reconfig_readdata[27]~9 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!Equal41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_reconfig_readdata[27]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_reconfig_readdata[27]~9 .extended_lut = "off";
defparam \user_reconfig_readdata[27]~9 .lut_mask = 64'h2028202820282028;
defparam \user_reconfig_readdata[27]~9 .shared_arith = "off";

dffeas \uif_writedata[25] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_25),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[25]~q ),
	.prn(vcc));
defparam \uif_writedata[25] .is_wysiwyg = "true";
defparam \uif_writedata[25] .power_up = "low";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\user_reconfig_readdata[27]~9_combout ),
	.datac(!\uif_writedata[25]~q ),
	.datad(!ph_readdata_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h0123012301230123;
defparam \Mux10~0 .shared_arith = "off";

dffeas \uif_writedata[26] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_26),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[26]~q ),
	.prn(vcc));
defparam \uif_writedata[26] .is_wysiwyg = "true";
defparam \uif_writedata[26] .power_up = "low";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\user_reconfig_readdata[27]~9_combout ),
	.datac(!\uif_writedata[26]~q ),
	.datad(!ph_readdata_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h0123012301230123;
defparam \Mux9~0 .shared_arith = "off";

dffeas \uif_writedata[27] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_27),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[27]~q ),
	.prn(vcc));
defparam \uif_writedata[27] .is_wysiwyg = "true";
defparam \uif_writedata[27] .power_up = "low";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\user_reconfig_readdata[27]~9_combout ),
	.datac(!\uif_writedata[27]~q ),
	.datad(!ph_readdata_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h0123012301230123;
defparam \Mux8~0 .shared_arith = "off";

dffeas \uif_writedata[28] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_28),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[28]~q ),
	.prn(vcc));
defparam \uif_writedata[28] .is_wysiwyg = "true";
defparam \uif_writedata[28] .power_up = "low";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\user_reconfig_readdata[27]~9_combout ),
	.datac(!\uif_writedata[28]~q ),
	.datad(!ph_readdata_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h0123012301230123;
defparam \Mux7~0 .shared_arith = "off";

dffeas \uif_writedata[29] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_29),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[29]~q ),
	.prn(vcc));
defparam \uif_writedata[29] .is_wysiwyg = "true";
defparam \uif_writedata[29] .power_up = "low";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\user_reconfig_readdata[27]~9_combout ),
	.datac(!\uif_writedata[29]~q ),
	.datad(!ph_readdata_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h0123012301230123;
defparam \Mux6~0 .shared_arith = "off";

dffeas \uif_writedata[30] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_30),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[30]~q ),
	.prn(vcc));
defparam \uif_writedata[30] .is_wysiwyg = "true";
defparam \uif_writedata[30] .power_up = "low";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\user_reconfig_readdata[27]~9_combout ),
	.datac(!\uif_writedata[30]~q ),
	.datad(!ph_readdata_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'h0123012301230123;
defparam \Mux5~0 .shared_arith = "off";

dffeas \uif_writedata[31] (
	.clk(mgmt_clk_clk),
	.d(reconfig_mgmt_writedata_31),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_writedata[0]~0_combout ),
	.q(\uif_writedata[31]~q ),
	.prn(vcc));
defparam \uif_writedata[31] .is_wysiwyg = "true";
defparam \uif_writedata[31] .power_up = "low";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!reconfig_mgmt_address_2),
	.datab(!\user_reconfig_readdata[27]~9_combout ),
	.datac(!\uif_writedata[31]~q ),
	.datad(!ph_readdata_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'h0123012301230123;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_mode[1]~1 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_mode[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_mode[1]~1 .extended_lut = "off";
defparam \uif_mode[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \uif_mode[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~1 (
	.dataa(!comb),
	.datab(!pll_mif_busy),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~1 .extended_lut = "off";
defparam \Mux0~1 .lut_mask = 64'h4444444444444444;
defparam \Mux0~1 .shared_arith = "off";

cyclonev_lcell_comb \uif_mode[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!uif_mode_01),
	.datac(!Mux0),
	.datad(!\always0~0_combout ),
	.datae(!\Mux0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_mode[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_mode[0]~0 .extended_lut = "off";
defparam \uif_mode[0]~0 .lut_mask = 64'h00040A0E00040A0E;
defparam \uif_mode[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_logical_ch_addr[0]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_logical_ch_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_logical_ch_addr[0]~0 .extended_lut = "off";
defparam \uif_logical_ch_addr[0]~0 .lut_mask = 64'h0080008000800080;
defparam \uif_logical_ch_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_addr_offset[2]~0 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!reconfig_mgmt_address_0),
	.datac(!reconfig_mgmt_address_2),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_addr_offset[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_addr_offset[2]~0 .extended_lut = "off";
defparam \uif_addr_offset[2]~0 .lut_mask = 64'h0010001000100010;
defparam \uif_addr_offset[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~2 (
	.dataa(!reconfig_mgmt_address_1),
	.datab(!uif_mode_01),
	.datac(!Mux0),
	.datad(!\always0~0_combout ),
	.datae(!\Mux0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~2 .extended_lut = "off";
defparam \Mux0~2 .lut_mask = 64'h00040A0E00040A0E;
defparam \Mux0~2 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_altera_wait_generate_3 (
	resync_chains0sync_r_1,
	launch_reg1,
	wait_reg1,
	ifsel_notdone_resync,
	launch_signal,
	mgmt_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
output 	launch_reg1;
output 	wait_reg1;
input 	ifsel_notdone_resync;
input 	launch_signal;
input 	mgmt_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_reg~0_combout ;


RECONFIGURE_IP_alt_xcvr_resync_3 rst_sync(
	.resync_chains0sync_r_1(resync_chains0sync_r_1),
	.ifsel_notdone_resync(ifsel_notdone_resync),
	.clk(mgmt_clk_clk));

dffeas launch_reg(
	.clk(mgmt_clk_clk),
	.d(launch_signal),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(launch_reg1),
	.prn(vcc));
defparam launch_reg.is_wysiwyg = "true";
defparam launch_reg.power_up = "low";

dffeas wait_reg(
	.clk(mgmt_clk_clk),
	.d(\wait_reg~0_combout ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_reg1),
	.prn(vcc));
defparam wait_reg.is_wysiwyg = "true";
defparam wait_reg.power_up = "low";

cyclonev_lcell_comb \wait_reg~0 (
	.dataa(!resync_chains0sync_r_1),
	.datab(!launch_signal),
	.datac(!launch_reg1),
	.datad(!wait_reg1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_reg~0 .extended_lut = "off";
defparam \wait_reg~0 .lut_mask = 64'h0100010001000100;
defparam \wait_reg~0 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_resync_3 (
	resync_chains0sync_r_1,
	ifsel_notdone_resync,
	clk)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
input 	ifsel_notdone_resync;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \resync_chains[0].sync_r[0]~q ;


dffeas \resync_chains[0].sync_r[1] (
	.clk(clk),
	.d(\resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resync_chains0sync_r_1),
	.prn(vcc));
defparam \resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[1] .power_up = "low";

dffeas \resync_chains[0].sync_r[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(ifsel_notdone_resync),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[0] .power_up = "low";

endmodule

module RECONFIGURE_IP_av_xcvr_reconfig_pll_ctrl (
	uif_rdata_3,
	uif_rdata_4,
	uif_rdata_5,
	uif_rdata_6,
	uif_rdata_7,
	uif_rdata_8,
	uif_rdata_9,
	uif_rdata_10,
	uif_rdata_11,
	uif_rdata_12,
	uif_rdata_13,
	uif_rdata_14,
	uif_rdata_15,
	uif_rdata_16,
	uif_rdata_17,
	uif_rdata_18,
	uif_rdata_19,
	ctrl_wdata_1,
	ctrl_addr_1,
	ctrl_wdata_2,
	ctrl_addr_5,
	ctrl_wdata_0,
	ctrl_addr_0,
	ctrl_addr_4,
	ctrl_wdata_5,
	ctrl_wdata_9,
	ctrl_wdata_13,
	ctrl_wdata_14,
	ctrl_wdata_15,
	pll_mif_busy1,
	reset,
	uif_logical_ch_addr_0,
	uif_wdata,
	uif_mode_1,
	uif_mode_0,
	Equal4,
	uif_rdata_0,
	uif_logical_ch_addr_01,
	uif_addr_offset_0,
	uif_logical_ch_addr_1,
	uif_rdata_1,
	uif_logical_ch_addr_11,
	uif_addr_offset_1,
	uif_logical_ch_addr_2,
	uif_rdata_2,
	uif_logical_ch_addr_21,
	uif_addr_offset_2,
	uif_logical_ch_addr_3,
	uif_logical_ch_addr_31,
	uif_logical_ch_addr_4,
	uif_logical_ch_addr_41,
	uif_logical_ch_addr_5,
	uif_logical_ch_addr_51,
	uif_logical_ch_addr_6,
	uif_logical_ch_addr_61,
	uif_logical_ch_addr_7,
	uif_logical_ch_addr_71,
	uif_logical_ch_addr_8,
	uif_logical_ch_addr_81,
	uif_logical_ch_addr_9,
	uif_logical_ch_addr_91,
	uif_addr_err1,
	uif_rdata_20,
	uif_rdata_21,
	uif_rdata_22,
	uif_rdata_23,
	uif_rdata_24,
	ctrl_go1,
	ctrl_lock1,
	ctrl_opcode_2,
	ctrl_opcode_0,
	pll_go,
	uif_go,
	waitrequest_to_ctrl,
	ctrl_lch_4,
	ctrl_lch_5,
	ctrl_lch_2,
	ctrl_lch_3,
	ctrl_lch_0,
	ctrl_lch_1,
	ctrl_lch_8,
	ctrl_lch_9,
	ctrl_lch_6,
	ctrl_lch_7,
	ctrl_wdata_3,
	ctrl_wdata_4,
	ctrl_wdata_6,
	ctrl_wdata_7,
	ctrl_wdata_8,
	ctrl_wdata_10,
	ctrl_wdata_11,
	ctrl_wdata_12,
	ctrl_rdata,
	pll_type,
	readdata_for_user_20,
	readdata_for_user_21,
	readdata_for_user_22,
	readdata_for_user_23,
	readdata_for_user_24,
	mif_rec_addr_7,
	mif_rec_addr_5,
	mif_rec_addr_6,
	clk)/* synthesis synthesis_greybox=0 */;
output 	uif_rdata_3;
output 	uif_rdata_4;
output 	uif_rdata_5;
output 	uif_rdata_6;
output 	uif_rdata_7;
output 	uif_rdata_8;
output 	uif_rdata_9;
output 	uif_rdata_10;
output 	uif_rdata_11;
output 	uif_rdata_12;
output 	uif_rdata_13;
output 	uif_rdata_14;
output 	uif_rdata_15;
output 	uif_rdata_16;
output 	uif_rdata_17;
output 	uif_rdata_18;
output 	uif_rdata_19;
output 	ctrl_wdata_1;
output 	ctrl_addr_1;
output 	ctrl_wdata_2;
output 	ctrl_addr_5;
output 	ctrl_wdata_0;
output 	ctrl_addr_0;
output 	ctrl_addr_4;
output 	ctrl_wdata_5;
output 	ctrl_wdata_9;
output 	ctrl_wdata_13;
output 	ctrl_wdata_14;
output 	ctrl_wdata_15;
output 	pll_mif_busy1;
input 	reset;
input 	uif_logical_ch_addr_0;
input 	[31:0] uif_wdata;
input 	uif_mode_1;
input 	uif_mode_0;
output 	Equal4;
output 	uif_rdata_0;
input 	uif_logical_ch_addr_01;
input 	uif_addr_offset_0;
input 	uif_logical_ch_addr_1;
output 	uif_rdata_1;
input 	uif_logical_ch_addr_11;
input 	uif_addr_offset_1;
input 	uif_logical_ch_addr_2;
output 	uif_rdata_2;
input 	uif_logical_ch_addr_21;
input 	uif_addr_offset_2;
input 	uif_logical_ch_addr_3;
input 	uif_logical_ch_addr_31;
input 	uif_logical_ch_addr_4;
input 	uif_logical_ch_addr_41;
input 	uif_logical_ch_addr_5;
input 	uif_logical_ch_addr_51;
input 	uif_logical_ch_addr_6;
input 	uif_logical_ch_addr_61;
input 	uif_logical_ch_addr_7;
input 	uif_logical_ch_addr_71;
input 	uif_logical_ch_addr_8;
input 	uif_logical_ch_addr_81;
input 	uif_logical_ch_addr_9;
input 	uif_logical_ch_addr_91;
output 	uif_addr_err1;
output 	uif_rdata_20;
output 	uif_rdata_21;
output 	uif_rdata_22;
output 	uif_rdata_23;
output 	uif_rdata_24;
output 	ctrl_go1;
output 	ctrl_lock1;
output 	ctrl_opcode_2;
output 	ctrl_opcode_0;
input 	pll_go;
input 	uif_go;
input 	waitrequest_to_ctrl;
output 	ctrl_lch_4;
output 	ctrl_lch_5;
output 	ctrl_lch_2;
output 	ctrl_lch_3;
output 	ctrl_lch_0;
output 	ctrl_lch_1;
output 	ctrl_lch_8;
output 	ctrl_lch_9;
output 	ctrl_lch_6;
output 	ctrl_lch_7;
output 	ctrl_wdata_3;
output 	ctrl_wdata_4;
output 	ctrl_wdata_6;
output 	ctrl_wdata_7;
output 	ctrl_wdata_8;
output 	ctrl_wdata_10;
output 	ctrl_wdata_11;
output 	ctrl_wdata_12;
input 	[31:0] ctrl_rdata;
input 	pll_type;
input 	readdata_for_user_20;
input 	readdata_for_user_21;
input 	readdata_for_user_22;
input 	readdata_for_user_23;
input 	readdata_for_user_24;
input 	mif_rec_addr_7;
input 	mif_rec_addr_5;
input 	mif_rec_addr_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal4~1_combout ;
wire \Equal3~0_combout ;
wire \always13~0_combout ;
wire \uif_l2p_active~0_combout ;
wire \uif_l2p_active~q ;
wire \state_event[0]~0_combout ;
wire \state_event[0]~1_combout ;
wire \state_event[2]~4_combout ;
wire \state_event[2]~q ;
wire \pll_next_state.PLL_WR~0_combout ;
wire \pll_next_state.PLL_WR~1_combout ;
wire \pll_state.PLL_WR~q ;
wire \uif_cgb_sel_wr~0_combout ;
wire \pll_uif_go~q ;
wire \pll_next_state.PLL_RD_L2P~0_combout ;
wire \pll_state.PLL_RD_L2P~q ;
wire \pll_next_state.PLL_RD~0_combout ;
wire \pll_state.PLL_RD~q ;
wire \ctrl_go~0_combout ;
wire \Selector2~0_combout ;
wire \pll_state.PLL_WAIT~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \pll_state.PLL_DECIDE~q ;
wire \state_event[0]~3_combout ;
wire \state_event[0]~q ;
wire \state_event[1]~2_combout ;
wire \state_event[1]~q ;
wire \pll_next_state.PLL_CHK_WORDS~0_combout ;
wire \pll_state.PLL_CHK_WORDS~q ;
wire \word_cnt~0_combout ;
wire \word_cnt[0]~q ;
wire \mif_req~0_combout ;
wire \mif_req~q ;
wire \pll_uif_type~0_combout ;
wire \pll_uif_type~1_combout ;
wire \pll_uif_type~q ;
wire \mux_pll_type~0_combout ;
wire \always6~0_combout ;
wire \phys_cgb[3]~q ;
wire \phys_refclk[0]~0_combout ;
wire \phys_refclk[3]~q ;
wire \phys_cgb[4]~q ;
wire \phys_refclk[4]~q ;
wire \phys_cgb[5]~q ;
wire \phys_refclk[5]~q ;
wire \phys_cgb[6]~q ;
wire \phys_refclk[6]~q ;
wire \phys_cgb[7]~q ;
wire \phys_refclk[7]~q ;
wire \phys_cgb[8]~q ;
wire \phys_refclk[8]~q ;
wire \phys_cgb[9]~q ;
wire \phys_refclk[9]~q ;
wire \phys_cgb[10]~q ;
wire \phys_refclk[10]~q ;
wire \phys_cgb[11]~q ;
wire \phys_refclk[11]~q ;
wire \phys_cgb[12]~q ;
wire \phys_refclk[12]~q ;
wire \phys_cgb[13]~q ;
wire \phys_refclk[13]~q ;
wire \phys_cgb[14]~q ;
wire \phys_refclk[14]~q ;
wire \phys_cgb[15]~q ;
wire \phys_refclk[15]~q ;
wire \phys_cgb[16]~q ;
wire \phys_refclk[16]~q ;
wire \phys_cgb[17]~q ;
wire \phys_refclk[17]~q ;
wire \phys_cgb[18]~q ;
wire \phys_refclk[18]~q ;
wire \phys_cgb[19]~q ;
wire \phys_refclk[19]~q ;
wire \modify_data[5]~0_combout ;
wire \phys_cgb[0]~q ;
wire \uif_rc_sel_wr~0_combout ;
wire \pll_uif_rc_sel[2]~q ;
wire \uif_cgb_sel_wr~1_combout ;
wire \pll_uif_cgb_sel[2]~q ;
wire \logical_index[2]~0_combout ;
wire \pll_uif_rc_sel[0]~q ;
wire \pll_uif_cgb_sel[0]~q ;
wire \logical_index[0]~1_combout ;
wire \pll_uif_rc_sel[1]~q ;
wire \pll_uif_cgb_sel[1]~q ;
wire \logical_index[1]~2_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux20~2_combout ;
wire \Mux21~2_combout ;
wire \phys_cgb[2]~q ;
wire \Mux21~3_combout ;
wire \Mux21~4_combout ;
wire \always11~0_combout ;
wire \saved_read_data[1]~q ;
wire \ctrl_wdata~0_combout ;
wire \ctrl_wdata[1]~1_combout ;
wire \ctrl_addr~0_combout ;
wire \ctrl_addr~1_combout ;
wire \Mux22~0_combout ;
wire \phys_cgb[1]~q ;
wire \Mux22~1_combout ;
wire \Mux22~2_combout ;
wire \saved_read_data[2]~q ;
wire \ctrl_wdata~24_combout ;
wire \ctrl_addr~2_combout ;
wire \ctrl_addr~3_combout ;
wire \saved_read_data[0]~q ;
wire \ctrl_wdata~2_combout ;
wire \ctrl_addr~4_combout ;
wire \ctrl_addr~5_combout ;
wire \WideOr1~0_combout ;
wire \saved_read_data[5]~q ;
wire \phys_refclk[2]~q ;
wire \phys_refclk[22]~q ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \phys_refclk[23]~q ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \phys_refclk[1]~q ;
wire \phys_refclk[21]~q ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \phys_refclk[0]~q ;
wire \phys_refclk[20]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \phys_refclk[24]~q ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \modify_data[5]~1_combout ;
wire \modify_data[5]~2_combout ;
wire \Ram0~3_combout ;
wire \saved_read_data[3]~q ;
wire \saved_read_data[9]~q ;
wire \WideOr0~0_combout ;
wire \modify_data[9]~3_combout ;
wire \saved_read_data[13]~q ;
wire \ctrl_wdata~17_combout ;
wire \saved_read_data[14]~q ;
wire \ctrl_wdata~18_combout ;
wire \saved_read_data[15]~q ;
wire \ctrl_wdata~19_combout ;
wire \Selector0~2_combout ;
wire \Selector0~3_combout ;
wire \Mux19~0_combout ;
wire \Mux18~0_combout ;
wire \Mux17~0_combout ;
wire \uif_rdata~0_combout ;
wire \uif_rdata~1_combout ;
wire \uif_rdata~2_combout ;
wire \uif_rdata~3_combout ;
wire \uif_rdata~4_combout ;
wire \ctrl_lock~0_combout ;
wire \ctrl_opcode[0]~0_combout ;
wire \ctrl_opcode~1_combout ;
wire \ctrl_wdata~3_combout ;
wire \ctrl_wdata[4]~4_combout ;
wire \ctrl_wdata[4]~5_combout ;
wire \WideOr2~0_combout ;
wire \ctrl_wdata~6_combout ;
wire \Ram0~0_combout ;
wire \saved_read_data[4]~q ;
wire \ctrl_wdata~7_combout ;
wire \ctrl_wdata~8_combout ;
wire \ctrl_wdata[6]~9_combout ;
wire \saved_read_data[6]~q ;
wire \ctrl_wdata~10_combout ;
wire \Ram0~1_combout ;
wire \saved_read_data[7]~q ;
wire \ctrl_wdata~11_combout ;
wire \Ram0~2_combout ;
wire \saved_read_data[8]~q ;
wire \ctrl_wdata~12_combout ;
wire \Ram0~4_combout ;
wire \saved_read_data[10]~q ;
wire \ctrl_wdata~13_combout ;
wire \ctrl_wdata~14_combout ;
wire \saved_read_data[11]~q ;
wire \ctrl_wdata~20_combout ;
wire \ctrl_wdata~15_combout ;
wire \saved_read_data[12]~q ;
wire \ctrl_wdata~16_combout ;


dffeas \uif_rdata[3] (
	.clk(clk),
	.d(\phys_cgb[3]~q ),
	.asdata(\phys_refclk[3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_3),
	.prn(vcc));
defparam \uif_rdata[3] .is_wysiwyg = "true";
defparam \uif_rdata[3] .power_up = "low";

dffeas \uif_rdata[4] (
	.clk(clk),
	.d(\phys_cgb[4]~q ),
	.asdata(\phys_refclk[4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_4),
	.prn(vcc));
defparam \uif_rdata[4] .is_wysiwyg = "true";
defparam \uif_rdata[4] .power_up = "low";

dffeas \uif_rdata[5] (
	.clk(clk),
	.d(\phys_cgb[5]~q ),
	.asdata(\phys_refclk[5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_5),
	.prn(vcc));
defparam \uif_rdata[5] .is_wysiwyg = "true";
defparam \uif_rdata[5] .power_up = "low";

dffeas \uif_rdata[6] (
	.clk(clk),
	.d(\phys_cgb[6]~q ),
	.asdata(\phys_refclk[6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_6),
	.prn(vcc));
defparam \uif_rdata[6] .is_wysiwyg = "true";
defparam \uif_rdata[6] .power_up = "low";

dffeas \uif_rdata[7] (
	.clk(clk),
	.d(\phys_cgb[7]~q ),
	.asdata(\phys_refclk[7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_7),
	.prn(vcc));
defparam \uif_rdata[7] .is_wysiwyg = "true";
defparam \uif_rdata[7] .power_up = "low";

dffeas \uif_rdata[8] (
	.clk(clk),
	.d(\phys_cgb[8]~q ),
	.asdata(\phys_refclk[8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_8),
	.prn(vcc));
defparam \uif_rdata[8] .is_wysiwyg = "true";
defparam \uif_rdata[8] .power_up = "low";

dffeas \uif_rdata[9] (
	.clk(clk),
	.d(\phys_cgb[9]~q ),
	.asdata(\phys_refclk[9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_9),
	.prn(vcc));
defparam \uif_rdata[9] .is_wysiwyg = "true";
defparam \uif_rdata[9] .power_up = "low";

dffeas \uif_rdata[10] (
	.clk(clk),
	.d(\phys_cgb[10]~q ),
	.asdata(\phys_refclk[10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_10),
	.prn(vcc));
defparam \uif_rdata[10] .is_wysiwyg = "true";
defparam \uif_rdata[10] .power_up = "low";

dffeas \uif_rdata[11] (
	.clk(clk),
	.d(\phys_cgb[11]~q ),
	.asdata(\phys_refclk[11]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_11),
	.prn(vcc));
defparam \uif_rdata[11] .is_wysiwyg = "true";
defparam \uif_rdata[11] .power_up = "low";

dffeas \uif_rdata[12] (
	.clk(clk),
	.d(\phys_cgb[12]~q ),
	.asdata(\phys_refclk[12]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_12),
	.prn(vcc));
defparam \uif_rdata[12] .is_wysiwyg = "true";
defparam \uif_rdata[12] .power_up = "low";

dffeas \uif_rdata[13] (
	.clk(clk),
	.d(\phys_cgb[13]~q ),
	.asdata(\phys_refclk[13]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_13),
	.prn(vcc));
defparam \uif_rdata[13] .is_wysiwyg = "true";
defparam \uif_rdata[13] .power_up = "low";

dffeas \uif_rdata[14] (
	.clk(clk),
	.d(\phys_cgb[14]~q ),
	.asdata(\phys_refclk[14]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_14),
	.prn(vcc));
defparam \uif_rdata[14] .is_wysiwyg = "true";
defparam \uif_rdata[14] .power_up = "low";

dffeas \uif_rdata[15] (
	.clk(clk),
	.d(\phys_cgb[15]~q ),
	.asdata(\phys_refclk[15]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_15),
	.prn(vcc));
defparam \uif_rdata[15] .is_wysiwyg = "true";
defparam \uif_rdata[15] .power_up = "low";

dffeas \uif_rdata[16] (
	.clk(clk),
	.d(\phys_cgb[16]~q ),
	.asdata(\phys_refclk[16]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_16),
	.prn(vcc));
defparam \uif_rdata[16] .is_wysiwyg = "true";
defparam \uif_rdata[16] .power_up = "low";

dffeas \uif_rdata[17] (
	.clk(clk),
	.d(\phys_cgb[17]~q ),
	.asdata(\phys_refclk[17]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_17),
	.prn(vcc));
defparam \uif_rdata[17] .is_wysiwyg = "true";
defparam \uif_rdata[17] .power_up = "low";

dffeas \uif_rdata[18] (
	.clk(clk),
	.d(\phys_cgb[18]~q ),
	.asdata(\phys_refclk[18]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_18),
	.prn(vcc));
defparam \uif_rdata[18] .is_wysiwyg = "true";
defparam \uif_rdata[18] .power_up = "low";

dffeas \uif_rdata[19] (
	.clk(clk),
	.d(\phys_cgb[19]~q ),
	.asdata(\phys_refclk[19]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal3~0_combout ),
	.sload(!uif_addr_offset_0),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_19),
	.prn(vcc));
defparam \uif_rdata[19] .is_wysiwyg = "true";
defparam \uif_rdata[19] .power_up = "low";

dffeas \ctrl_wdata[1] (
	.clk(clk),
	.d(\ctrl_wdata~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_1),
	.prn(vcc));
defparam \ctrl_wdata[1] .is_wysiwyg = "true";
defparam \ctrl_wdata[1] .power_up = "low";

dffeas \ctrl_addr[1] (
	.clk(clk),
	.d(\ctrl_addr~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_addr~1_combout ),
	.q(ctrl_addr_1),
	.prn(vcc));
defparam \ctrl_addr[1] .is_wysiwyg = "true";
defparam \ctrl_addr[1] .power_up = "low";

dffeas \ctrl_wdata[2] (
	.clk(clk),
	.d(\ctrl_wdata~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_2),
	.prn(vcc));
defparam \ctrl_wdata[2] .is_wysiwyg = "true";
defparam \ctrl_wdata[2] .power_up = "low";

dffeas \ctrl_addr[5] (
	.clk(clk),
	.d(\ctrl_addr~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_addr~1_combout ),
	.q(ctrl_addr_5),
	.prn(vcc));
defparam \ctrl_addr[5] .is_wysiwyg = "true";
defparam \ctrl_addr[5] .power_up = "low";

dffeas \ctrl_wdata[0] (
	.clk(clk),
	.d(\ctrl_wdata~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_0),
	.prn(vcc));
defparam \ctrl_wdata[0] .is_wysiwyg = "true";
defparam \ctrl_wdata[0] .power_up = "low";

dffeas \ctrl_addr[0] (
	.clk(clk),
	.d(\ctrl_addr~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_addr~1_combout ),
	.q(ctrl_addr_0),
	.prn(vcc));
defparam \ctrl_addr[0] .is_wysiwyg = "true";
defparam \ctrl_addr[0] .power_up = "low";

dffeas \ctrl_addr[4] (
	.clk(clk),
	.d(\ctrl_addr~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_addr~1_combout ),
	.q(ctrl_addr_4),
	.prn(vcc));
defparam \ctrl_addr[4] .is_wysiwyg = "true";
defparam \ctrl_addr[4] .power_up = "low";

dffeas \ctrl_wdata[5] (
	.clk(clk),
	.d(\modify_data[5]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_5),
	.prn(vcc));
defparam \ctrl_wdata[5] .is_wysiwyg = "true";
defparam \ctrl_wdata[5] .power_up = "low";

dffeas \ctrl_wdata[9] (
	.clk(clk),
	.d(\modify_data[9]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_9),
	.prn(vcc));
defparam \ctrl_wdata[9] .is_wysiwyg = "true";
defparam \ctrl_wdata[9] .power_up = "low";

dffeas \ctrl_wdata[13] (
	.clk(clk),
	.d(\ctrl_wdata~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_13),
	.prn(vcc));
defparam \ctrl_wdata[13] .is_wysiwyg = "true";
defparam \ctrl_wdata[13] .power_up = "low";

dffeas \ctrl_wdata[14] (
	.clk(clk),
	.d(\ctrl_wdata~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_14),
	.prn(vcc));
defparam \ctrl_wdata[14] .is_wysiwyg = "true";
defparam \ctrl_wdata[14] .power_up = "low";

dffeas \ctrl_wdata[15] (
	.clk(clk),
	.d(\ctrl_wdata~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!pll_mif_busy1),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_15),
	.prn(vcc));
defparam \ctrl_wdata[15] .is_wysiwyg = "true";
defparam \ctrl_wdata[15] .power_up = "low";

dffeas pll_mif_busy(
	.clk(clk),
	.d(\Selector0~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pll_mif_busy1),
	.prn(vcc));
defparam pll_mif_busy.is_wysiwyg = "true";
defparam pll_mif_busy.power_up = "low";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h2222222222222222;
defparam \Equal4~0 .shared_arith = "off";

dffeas \uif_rdata[0] (
	.clk(clk),
	.d(\Mux19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_0),
	.prn(vcc));
defparam \uif_rdata[0] .is_wysiwyg = "true";
defparam \uif_rdata[0] .power_up = "low";

dffeas \uif_rdata[1] (
	.clk(clk),
	.d(\Mux18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_1),
	.prn(vcc));
defparam \uif_rdata[1] .is_wysiwyg = "true";
defparam \uif_rdata[1] .power_up = "low";

dffeas \uif_rdata[2] (
	.clk(clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_2),
	.prn(vcc));
defparam \uif_rdata[2] .is_wysiwyg = "true";
defparam \uif_rdata[2] .power_up = "low";

dffeas uif_addr_err(
	.clk(clk),
	.d(uif_addr_offset_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(uif_addr_err1),
	.prn(vcc));
defparam uif_addr_err.is_wysiwyg = "true";
defparam uif_addr_err.power_up = "low";

dffeas \uif_rdata[20] (
	.clk(clk),
	.d(\uif_rdata~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_20),
	.prn(vcc));
defparam \uif_rdata[20] .is_wysiwyg = "true";
defparam \uif_rdata[20] .power_up = "low";

dffeas \uif_rdata[21] (
	.clk(clk),
	.d(\uif_rdata~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_21),
	.prn(vcc));
defparam \uif_rdata[21] .is_wysiwyg = "true";
defparam \uif_rdata[21] .power_up = "low";

dffeas \uif_rdata[22] (
	.clk(clk),
	.d(\uif_rdata~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_22),
	.prn(vcc));
defparam \uif_rdata[22] .is_wysiwyg = "true";
defparam \uif_rdata[22] .power_up = "low";

dffeas \uif_rdata[23] (
	.clk(clk),
	.d(\uif_rdata~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_23),
	.prn(vcc));
defparam \uif_rdata[23] .is_wysiwyg = "true";
defparam \uif_rdata[23] .power_up = "low";

dffeas \uif_rdata[24] (
	.clk(clk),
	.d(\uif_rdata~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal4~1_combout ),
	.q(uif_rdata_24),
	.prn(vcc));
defparam \uif_rdata[24] .is_wysiwyg = "true";
defparam \uif_rdata[24] .power_up = "low";

dffeas ctrl_go(
	.clk(clk),
	.d(\ctrl_go~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_go1),
	.prn(vcc));
defparam ctrl_go.is_wysiwyg = "true";
defparam ctrl_go.power_up = "low";

dffeas ctrl_lock(
	.clk(clk),
	.d(\ctrl_lock~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctrl_lock1),
	.prn(vcc));
defparam ctrl_lock.is_wysiwyg = "true";
defparam ctrl_lock.power_up = "low";

dffeas \ctrl_opcode[2] (
	.clk(clk),
	.d(\pll_state.PLL_RD_L2P~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_opcode[0]~0_combout ),
	.q(ctrl_opcode_2),
	.prn(vcc));
defparam \ctrl_opcode[2] .is_wysiwyg = "true";
defparam \ctrl_opcode[2] .power_up = "low";

dffeas \ctrl_opcode[0] (
	.clk(clk),
	.d(\ctrl_opcode~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_opcode[0]~0_combout ),
	.q(ctrl_opcode_0),
	.prn(vcc));
defparam \ctrl_opcode[0] .is_wysiwyg = "true";
defparam \ctrl_opcode[0] .power_up = "low";

cyclonev_lcell_comb \ctrl_lch[4]~0 (
	.dataa(!uif_logical_ch_addr_4),
	.datab(!uif_logical_ch_addr_41),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[4]~0 .extended_lut = "off";
defparam \ctrl_lch[4]~0 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[5]~1 (
	.dataa(!uif_logical_ch_addr_5),
	.datab(!uif_logical_ch_addr_51),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[5]~1 .extended_lut = "off";
defparam \ctrl_lch[5]~1 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[2]~2 (
	.dataa(!uif_logical_ch_addr_2),
	.datab(!uif_logical_ch_addr_21),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[2]~2 .extended_lut = "off";
defparam \ctrl_lch[2]~2 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[3]~3 (
	.dataa(!uif_logical_ch_addr_3),
	.datab(!uif_logical_ch_addr_31),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[3]~3 .extended_lut = "off";
defparam \ctrl_lch[3]~3 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[0]~4 (
	.dataa(!uif_logical_ch_addr_0),
	.datab(!uif_logical_ch_addr_01),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[0]~4 .extended_lut = "off";
defparam \ctrl_lch[0]~4 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[1]~5 (
	.dataa(!uif_logical_ch_addr_1),
	.datab(!uif_logical_ch_addr_11),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[1]~5 .extended_lut = "off";
defparam \ctrl_lch[1]~5 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[1]~5 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[8]~6 (
	.dataa(!uif_logical_ch_addr_81),
	.datab(!uif_logical_ch_addr_8),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[8]~6 .extended_lut = "off";
defparam \ctrl_lch[8]~6 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[8]~6 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[9]~7 (
	.dataa(!uif_logical_ch_addr_9),
	.datab(!uif_logical_ch_addr_91),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[9]~7 .extended_lut = "off";
defparam \ctrl_lch[9]~7 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[9]~7 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[6]~8 (
	.dataa(!uif_logical_ch_addr_6),
	.datab(!uif_logical_ch_addr_61),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[6]~8 .extended_lut = "off";
defparam \ctrl_lch[6]~8 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lch[7]~9 (
	.dataa(!uif_logical_ch_addr_7),
	.datab(!uif_logical_ch_addr_71),
	.datac(!\mif_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_lch_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lch[7]~9 .extended_lut = "off";
defparam \ctrl_lch[7]~9 .lut_mask = 64'h3535353535353535;
defparam \ctrl_lch[7]~9 .shared_arith = "off";

dffeas \ctrl_wdata[3] (
	.clk(clk),
	.d(\ctrl_wdata~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_3),
	.prn(vcc));
defparam \ctrl_wdata[3] .is_wysiwyg = "true";
defparam \ctrl_wdata[3] .power_up = "low";

dffeas \ctrl_wdata[4] (
	.clk(clk),
	.d(\ctrl_wdata~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_4),
	.prn(vcc));
defparam \ctrl_wdata[4] .is_wysiwyg = "true";
defparam \ctrl_wdata[4] .power_up = "low";

dffeas \ctrl_wdata[6] (
	.clk(clk),
	.d(\ctrl_wdata~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_6),
	.prn(vcc));
defparam \ctrl_wdata[6] .is_wysiwyg = "true";
defparam \ctrl_wdata[6] .power_up = "low";

dffeas \ctrl_wdata[7] (
	.clk(clk),
	.d(\ctrl_wdata~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_7),
	.prn(vcc));
defparam \ctrl_wdata[7] .is_wysiwyg = "true";
defparam \ctrl_wdata[7] .power_up = "low";

dffeas \ctrl_wdata[8] (
	.clk(clk),
	.d(\ctrl_wdata~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_8),
	.prn(vcc));
defparam \ctrl_wdata[8] .is_wysiwyg = "true";
defparam \ctrl_wdata[8] .power_up = "low";

dffeas \ctrl_wdata[10] (
	.clk(clk),
	.d(\ctrl_wdata~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_10),
	.prn(vcc));
defparam \ctrl_wdata[10] .is_wysiwyg = "true";
defparam \ctrl_wdata[10] .power_up = "low";

dffeas \ctrl_wdata[11] (
	.clk(clk),
	.d(\ctrl_wdata~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_11),
	.prn(vcc));
defparam \ctrl_wdata[11] .is_wysiwyg = "true";
defparam \ctrl_wdata[11] .power_up = "low";

dffeas \ctrl_wdata[12] (
	.clk(clk),
	.d(\ctrl_wdata~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ctrl_wdata[1]~1_combout ),
	.q(ctrl_wdata_12),
	.prn(vcc));
defparam \ctrl_wdata[12] .is_wysiwyg = "true";
defparam \ctrl_wdata[12] .power_up = "low";

cyclonev_lcell_comb \Equal4~1 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'h8888888888888888;
defparam \Equal4~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!uif_addr_offset_1),
	.datab(!uif_addr_offset_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \always13~0 (
	.dataa(!uif_go),
	.datab(!\Equal4~1_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~0 .extended_lut = "off";
defparam \always13~0 .lut_mask = 64'h1010101010101010;
defparam \always13~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_l2p_active~0 (
	.dataa(!\always13~0_combout ),
	.datab(!\uif_l2p_active~q ),
	.datac(!waitrequest_to_ctrl),
	.datad(!\pll_state.PLL_DECIDE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_l2p_active~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_l2p_active~0 .extended_lut = "off";
defparam \uif_l2p_active~0 .lut_mask = 64'h7747774777477747;
defparam \uif_l2p_active~0 .shared_arith = "off";

dffeas uif_l2p_active(
	.clk(clk),
	.d(\uif_l2p_active~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\uif_l2p_active~q ),
	.prn(vcc));
defparam uif_l2p_active.is_wysiwyg = "true";
defparam uif_l2p_active.power_up = "low";

cyclonev_lcell_comb \state_event[0]~0 (
	.dataa(!\uif_l2p_active~q ),
	.datab(!waitrequest_to_ctrl),
	.datac(!\state_event[1]~q ),
	.datad(!\state_event[0]~q ),
	.datae(!\state_event[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state_event[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state_event[0]~0 .extended_lut = "off";
defparam \state_event[0]~0 .lut_mask = 64'h0008000000080000;
defparam \state_event[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \state_event[0]~1 (
	.dataa(!pll_mif_busy1),
	.datab(!\pll_state.PLL_DECIDE~q ),
	.datac(!\pll_state.PLL_WAIT~q ),
	.datad(!\state_event[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state_event[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state_event[0]~1 .extended_lut = "off";
defparam \state_event[0]~1 .lut_mask = 64'h5140514051405140;
defparam \state_event[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \state_event[2]~4 (
	.dataa(!pll_mif_busy1),
	.datab(!\state_event[1]~q ),
	.datac(!\state_event[0]~q ),
	.datad(!\state_event[2]~q ),
	.datae(!\pll_next_state.PLL_WR~0_combout ),
	.dataf(!\state_event[0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state_event[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state_event[2]~4 .extended_lut = "off";
defparam \state_event[2]~4 .lut_mask = 64'h0154005400FF00FF;
defparam \state_event[2]~4 .shared_arith = "off";

dffeas \state_event[2] (
	.clk(clk),
	.d(\state_event[2]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_event[2]~q ),
	.prn(vcc));
defparam \state_event[2] .is_wysiwyg = "true";
defparam \state_event[2] .power_up = "low";

cyclonev_lcell_comb \pll_next_state.PLL_WR~0 (
	.dataa(!\uif_l2p_active~q ),
	.datab(!waitrequest_to_ctrl),
	.datac(!\pll_state.PLL_DECIDE~q ),
	.datad(!\state_event[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_next_state.PLL_WR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_next_state.PLL_WR~0 .extended_lut = "off";
defparam \pll_next_state.PLL_WR~0 .lut_mask = 64'h0800080008000800;
defparam \pll_next_state.PLL_WR~0 .shared_arith = "off";

cyclonev_lcell_comb \pll_next_state.PLL_WR~1 (
	.dataa(!\state_event[1]~q ),
	.datab(!\state_event[0]~q ),
	.datac(!\pll_next_state.PLL_WR~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_next_state.PLL_WR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_next_state.PLL_WR~1 .extended_lut = "off";
defparam \pll_next_state.PLL_WR~1 .lut_mask = 64'h0404040404040404;
defparam \pll_next_state.PLL_WR~1 .shared_arith = "off";

dffeas \pll_state.PLL_WR (
	.clk(clk),
	.d(\pll_next_state.PLL_WR~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_state.PLL_WR~q ),
	.prn(vcc));
defparam \pll_state.PLL_WR .is_wysiwyg = "true";
defparam \pll_state.PLL_WR .power_up = "low";

cyclonev_lcell_comb \uif_cgb_sel_wr~0 (
	.dataa(!Equal4),
	.datab(!uif_addr_offset_1),
	.datac(!uif_addr_offset_2),
	.datad(!uif_go),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_cgb_sel_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_cgb_sel_wr~0 .extended_lut = "off";
defparam \uif_cgb_sel_wr~0 .lut_mask = 64'h0040004000400040;
defparam \uif_cgb_sel_wr~0 .shared_arith = "off";

dffeas pll_uif_go(
	.clk(clk),
	.d(\uif_cgb_sel_wr~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_uif_go~q ),
	.prn(vcc));
defparam pll_uif_go.is_wysiwyg = "true";
defparam pll_uif_go.power_up = "low";

cyclonev_lcell_comb \pll_next_state.PLL_RD_L2P~0 (
	.dataa(!pll_mif_busy1),
	.datab(!pll_go),
	.datac(!\pll_uif_go~q ),
	.datad(!\always13~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_next_state.PLL_RD_L2P~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_next_state.PLL_RD_L2P~0 .extended_lut = "off";
defparam \pll_next_state.PLL_RD_L2P~0 .lut_mask = 64'h2AAA2AAA2AAA2AAA;
defparam \pll_next_state.PLL_RD_L2P~0 .shared_arith = "off";

dffeas \pll_state.PLL_RD_L2P (
	.clk(clk),
	.d(\pll_next_state.PLL_RD_L2P~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_state.PLL_RD_L2P~q ),
	.prn(vcc));
defparam \pll_state.PLL_RD_L2P .is_wysiwyg = "true";
defparam \pll_state.PLL_RD_L2P .power_up = "low";

cyclonev_lcell_comb \pll_next_state.PLL_RD~0 (
	.dataa(!\state_event[1]~q ),
	.datab(!\state_event[0]~q ),
	.datac(!\pll_next_state.PLL_WR~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_next_state.PLL_RD~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_next_state.PLL_RD~0 .extended_lut = "off";
defparam \pll_next_state.PLL_RD~0 .lut_mask = 64'h0202020202020202;
defparam \pll_next_state.PLL_RD~0 .shared_arith = "off";

dffeas \pll_state.PLL_RD (
	.clk(clk),
	.d(\pll_next_state.PLL_RD~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_state.PLL_RD~q ),
	.prn(vcc));
defparam \pll_state.PLL_RD .is_wysiwyg = "true";
defparam \pll_state.PLL_RD .power_up = "low";

cyclonev_lcell_comb \ctrl_go~0 (
	.dataa(!\pll_state.PLL_WR~q ),
	.datab(!\pll_state.PLL_RD_L2P~q ),
	.datac(!\pll_state.PLL_RD~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_go~0 .extended_lut = "off";
defparam \ctrl_go~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ctrl_go~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\pll_state.PLL_CHK_WORDS~q ),
	.datac(!\ctrl_go~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \Selector2~0 .shared_arith = "off";

dffeas \pll_state.PLL_WAIT (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_state.PLL_WAIT~q ),
	.prn(vcc));
defparam \pll_state.PLL_WAIT .is_wysiwyg = "true";
defparam \pll_state.PLL_WAIT .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\uif_l2p_active~q ),
	.datab(!\state_event[1]~q ),
	.datac(!\state_event[0]~q ),
	.datad(!\state_event[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h80AA80AA80AA80AA;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!waitrequest_to_ctrl),
	.datab(!\pll_state.PLL_DECIDE~q ),
	.datac(!\pll_state.PLL_WAIT~q ),
	.datad(!\Selector1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h1F3F1F3F1F3F1F3F;
defparam \Selector1~1 .shared_arith = "off";

dffeas \pll_state.PLL_DECIDE (
	.clk(clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_state.PLL_DECIDE~q ),
	.prn(vcc));
defparam \pll_state.PLL_DECIDE .is_wysiwyg = "true";
defparam \pll_state.PLL_DECIDE .power_up = "low";

cyclonev_lcell_comb \state_event[0]~3 (
	.dataa(!pll_mif_busy1),
	.datab(!\pll_state.PLL_DECIDE~q ),
	.datac(!\state_event[0]~q ),
	.datad(!\pll_state.PLL_WAIT~q ),
	.datae(!\state_event[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state_event[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state_event[0]~3 .extended_lut = "off";
defparam \state_event[0]~3 .lut_mask = 64'h0541044005410440;
defparam \state_event[0]~3 .shared_arith = "off";

dffeas \state_event[0] (
	.clk(clk),
	.d(\state_event[0]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_event[0]~q ),
	.prn(vcc));
defparam \state_event[0] .is_wysiwyg = "true";
defparam \state_event[0] .power_up = "low";

cyclonev_lcell_comb \state_event[1]~2 (
	.dataa(!pll_mif_busy1),
	.datab(!\state_event[1]~q ),
	.datac(!\state_event[0]~q ),
	.datad(gnd),
	.datae(!\state_event[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state_event[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state_event[1]~2 .extended_lut = "off";
defparam \state_event[1]~2 .lut_mask = 64'h1414333314143333;
defparam \state_event[1]~2 .shared_arith = "off";

dffeas \state_event[1] (
	.clk(clk),
	.d(\state_event[1]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_event[1]~q ),
	.prn(vcc));
defparam \state_event[1] .is_wysiwyg = "true";
defparam \state_event[1] .power_up = "low";

cyclonev_lcell_comb \pll_next_state.PLL_CHK_WORDS~0 (
	.dataa(!\state_event[1]~q ),
	.datab(!\state_event[0]~q ),
	.datac(!\pll_next_state.PLL_WR~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_next_state.PLL_CHK_WORDS~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_next_state.PLL_CHK_WORDS~0 .extended_lut = "off";
defparam \pll_next_state.PLL_CHK_WORDS~0 .lut_mask = 64'h0101010101010101;
defparam \pll_next_state.PLL_CHK_WORDS~0 .shared_arith = "off";

dffeas \pll_state.PLL_CHK_WORDS (
	.clk(clk),
	.d(\pll_next_state.PLL_CHK_WORDS~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_state.PLL_CHK_WORDS~q ),
	.prn(vcc));
defparam \pll_state.PLL_CHK_WORDS .is_wysiwyg = "true";
defparam \pll_state.PLL_CHK_WORDS .power_up = "low";

cyclonev_lcell_comb \word_cnt~0 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\pll_state.PLL_CHK_WORDS~q ),
	.datac(!\pll_state.PLL_RD_L2P~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\word_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \word_cnt~0 .extended_lut = "off";
defparam \word_cnt~0 .lut_mask = 64'h4F4F4F4F4F4F4F4F;
defparam \word_cnt~0 .shared_arith = "off";

dffeas \word_cnt[0] (
	.clk(clk),
	.d(\word_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\word_cnt[0]~q ),
	.prn(vcc));
defparam \word_cnt[0] .is_wysiwyg = "true";
defparam \word_cnt[0] .power_up = "low";

cyclonev_lcell_comb \mif_req~0 (
	.dataa(!pll_go),
	.datab(!\word_cnt[0]~q ),
	.datac(!\pll_state.PLL_CHK_WORDS~q ),
	.datad(!\mif_req~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mif_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mif_req~0 .extended_lut = "off";
defparam \mif_req~0 .lut_mask = 64'h51F351F351F351F3;
defparam \mif_req~0 .shared_arith = "off";

dffeas mif_req(
	.clk(clk),
	.d(\mif_req~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mif_req~q ),
	.prn(vcc));
defparam mif_req.is_wysiwyg = "true";
defparam mif_req.power_up = "low";

cyclonev_lcell_comb \pll_uif_type~0 (
	.dataa(!uif_mode_1),
	.datab(!uif_mode_0),
	.datac(!uif_addr_offset_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_uif_type~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_uif_type~0 .extended_lut = "off";
defparam \pll_uif_type~0 .lut_mask = 64'h2828282828282828;
defparam \pll_uif_type~0 .shared_arith = "off";

cyclonev_lcell_comb \pll_uif_type~1 (
	.dataa(!uif_addr_offset_0),
	.datab(!uif_addr_offset_2),
	.datac(!uif_go),
	.datad(!\pll_uif_type~q ),
	.datae(!\pll_uif_type~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_uif_type~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_uif_type~1 .extended_lut = "off";
defparam \pll_uif_type~1 .lut_mask = 64'h00FF04F700FF04F7;
defparam \pll_uif_type~1 .shared_arith = "off";

dffeas pll_uif_type(
	.clk(clk),
	.d(\pll_uif_type~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_uif_type~q ),
	.prn(vcc));
defparam pll_uif_type.is_wysiwyg = "true";
defparam pll_uif_type.power_up = "low";

cyclonev_lcell_comb \mux_pll_type~0 (
	.dataa(!\mif_req~q ),
	.datab(!pll_type),
	.datac(!\pll_uif_type~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mux_pll_type~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mux_pll_type~0 .extended_lut = "off";
defparam \mux_pll_type~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mux_pll_type~0 .shared_arith = "off";

cyclonev_lcell_comb \always6~0 (
	.dataa(!ctrl_opcode_2),
	.datab(!ctrl_opcode_0),
	.datac(!waitrequest_to_ctrl),
	.datad(!\mux_pll_type~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'h0040004000400040;
defparam \always6~0 .shared_arith = "off";

dffeas \phys_cgb[3] (
	.clk(clk),
	.d(ctrl_rdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[3]~q ),
	.prn(vcc));
defparam \phys_cgb[3] .is_wysiwyg = "true";
defparam \phys_cgb[3] .power_up = "low";

cyclonev_lcell_comb \phys_refclk[0]~0 (
	.dataa(!ctrl_opcode_2),
	.datab(!ctrl_opcode_0),
	.datac(!waitrequest_to_ctrl),
	.datad(!\mux_pll_type~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\phys_refclk[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \phys_refclk[0]~0 .extended_lut = "off";
defparam \phys_refclk[0]~0 .lut_mask = 64'h4000400040004000;
defparam \phys_refclk[0]~0 .shared_arith = "off";

dffeas \phys_refclk[3] (
	.clk(clk),
	.d(ctrl_rdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[3]~q ),
	.prn(vcc));
defparam \phys_refclk[3] .is_wysiwyg = "true";
defparam \phys_refclk[3] .power_up = "low";

dffeas \phys_cgb[4] (
	.clk(clk),
	.d(ctrl_rdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[4]~q ),
	.prn(vcc));
defparam \phys_cgb[4] .is_wysiwyg = "true";
defparam \phys_cgb[4] .power_up = "low";

dffeas \phys_refclk[4] (
	.clk(clk),
	.d(ctrl_rdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[4]~q ),
	.prn(vcc));
defparam \phys_refclk[4] .is_wysiwyg = "true";
defparam \phys_refclk[4] .power_up = "low";

dffeas \phys_cgb[5] (
	.clk(clk),
	.d(ctrl_rdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[5]~q ),
	.prn(vcc));
defparam \phys_cgb[5] .is_wysiwyg = "true";
defparam \phys_cgb[5] .power_up = "low";

dffeas \phys_refclk[5] (
	.clk(clk),
	.d(ctrl_rdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[5]~q ),
	.prn(vcc));
defparam \phys_refclk[5] .is_wysiwyg = "true";
defparam \phys_refclk[5] .power_up = "low";

dffeas \phys_cgb[6] (
	.clk(clk),
	.d(ctrl_rdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[6]~q ),
	.prn(vcc));
defparam \phys_cgb[6] .is_wysiwyg = "true";
defparam \phys_cgb[6] .power_up = "low";

dffeas \phys_refclk[6] (
	.clk(clk),
	.d(ctrl_rdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[6]~q ),
	.prn(vcc));
defparam \phys_refclk[6] .is_wysiwyg = "true";
defparam \phys_refclk[6] .power_up = "low";

dffeas \phys_cgb[7] (
	.clk(clk),
	.d(ctrl_rdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[7]~q ),
	.prn(vcc));
defparam \phys_cgb[7] .is_wysiwyg = "true";
defparam \phys_cgb[7] .power_up = "low";

dffeas \phys_refclk[7] (
	.clk(clk),
	.d(ctrl_rdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[7]~q ),
	.prn(vcc));
defparam \phys_refclk[7] .is_wysiwyg = "true";
defparam \phys_refclk[7] .power_up = "low";

dffeas \phys_cgb[8] (
	.clk(clk),
	.d(ctrl_rdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[8]~q ),
	.prn(vcc));
defparam \phys_cgb[8] .is_wysiwyg = "true";
defparam \phys_cgb[8] .power_up = "low";

dffeas \phys_refclk[8] (
	.clk(clk),
	.d(ctrl_rdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[8]~q ),
	.prn(vcc));
defparam \phys_refclk[8] .is_wysiwyg = "true";
defparam \phys_refclk[8] .power_up = "low";

dffeas \phys_cgb[9] (
	.clk(clk),
	.d(ctrl_rdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[9]~q ),
	.prn(vcc));
defparam \phys_cgb[9] .is_wysiwyg = "true";
defparam \phys_cgb[9] .power_up = "low";

dffeas \phys_refclk[9] (
	.clk(clk),
	.d(ctrl_rdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[9]~q ),
	.prn(vcc));
defparam \phys_refclk[9] .is_wysiwyg = "true";
defparam \phys_refclk[9] .power_up = "low";

dffeas \phys_cgb[10] (
	.clk(clk),
	.d(ctrl_rdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[10]~q ),
	.prn(vcc));
defparam \phys_cgb[10] .is_wysiwyg = "true";
defparam \phys_cgb[10] .power_up = "low";

dffeas \phys_refclk[10] (
	.clk(clk),
	.d(ctrl_rdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[10]~q ),
	.prn(vcc));
defparam \phys_refclk[10] .is_wysiwyg = "true";
defparam \phys_refclk[10] .power_up = "low";

dffeas \phys_cgb[11] (
	.clk(clk),
	.d(ctrl_rdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[11]~q ),
	.prn(vcc));
defparam \phys_cgb[11] .is_wysiwyg = "true";
defparam \phys_cgb[11] .power_up = "low";

dffeas \phys_refclk[11] (
	.clk(clk),
	.d(ctrl_rdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[11]~q ),
	.prn(vcc));
defparam \phys_refclk[11] .is_wysiwyg = "true";
defparam \phys_refclk[11] .power_up = "low";

dffeas \phys_cgb[12] (
	.clk(clk),
	.d(ctrl_rdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[12]~q ),
	.prn(vcc));
defparam \phys_cgb[12] .is_wysiwyg = "true";
defparam \phys_cgb[12] .power_up = "low";

dffeas \phys_refclk[12] (
	.clk(clk),
	.d(ctrl_rdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[12]~q ),
	.prn(vcc));
defparam \phys_refclk[12] .is_wysiwyg = "true";
defparam \phys_refclk[12] .power_up = "low";

dffeas \phys_cgb[13] (
	.clk(clk),
	.d(ctrl_rdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[13]~q ),
	.prn(vcc));
defparam \phys_cgb[13] .is_wysiwyg = "true";
defparam \phys_cgb[13] .power_up = "low";

dffeas \phys_refclk[13] (
	.clk(clk),
	.d(ctrl_rdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[13]~q ),
	.prn(vcc));
defparam \phys_refclk[13] .is_wysiwyg = "true";
defparam \phys_refclk[13] .power_up = "low";

dffeas \phys_cgb[14] (
	.clk(clk),
	.d(ctrl_rdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[14]~q ),
	.prn(vcc));
defparam \phys_cgb[14] .is_wysiwyg = "true";
defparam \phys_cgb[14] .power_up = "low";

dffeas \phys_refclk[14] (
	.clk(clk),
	.d(ctrl_rdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[14]~q ),
	.prn(vcc));
defparam \phys_refclk[14] .is_wysiwyg = "true";
defparam \phys_refclk[14] .power_up = "low";

dffeas \phys_cgb[15] (
	.clk(clk),
	.d(ctrl_rdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[15]~q ),
	.prn(vcc));
defparam \phys_cgb[15] .is_wysiwyg = "true";
defparam \phys_cgb[15] .power_up = "low";

dffeas \phys_refclk[15] (
	.clk(clk),
	.d(ctrl_rdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[15]~q ),
	.prn(vcc));
defparam \phys_refclk[15] .is_wysiwyg = "true";
defparam \phys_refclk[15] .power_up = "low";

dffeas \phys_cgb[16] (
	.clk(clk),
	.d(ctrl_rdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[16]~q ),
	.prn(vcc));
defparam \phys_cgb[16] .is_wysiwyg = "true";
defparam \phys_cgb[16] .power_up = "low";

dffeas \phys_refclk[16] (
	.clk(clk),
	.d(ctrl_rdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[16]~q ),
	.prn(vcc));
defparam \phys_refclk[16] .is_wysiwyg = "true";
defparam \phys_refclk[16] .power_up = "low";

dffeas \phys_cgb[17] (
	.clk(clk),
	.d(ctrl_rdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[17]~q ),
	.prn(vcc));
defparam \phys_cgb[17] .is_wysiwyg = "true";
defparam \phys_cgb[17] .power_up = "low";

dffeas \phys_refclk[17] (
	.clk(clk),
	.d(ctrl_rdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[17]~q ),
	.prn(vcc));
defparam \phys_refclk[17] .is_wysiwyg = "true";
defparam \phys_refclk[17] .power_up = "low";

dffeas \phys_cgb[18] (
	.clk(clk),
	.d(ctrl_rdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[18]~q ),
	.prn(vcc));
defparam \phys_cgb[18] .is_wysiwyg = "true";
defparam \phys_cgb[18] .power_up = "low";

dffeas \phys_refclk[18] (
	.clk(clk),
	.d(ctrl_rdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[18]~q ),
	.prn(vcc));
defparam \phys_refclk[18] .is_wysiwyg = "true";
defparam \phys_refclk[18] .power_up = "low";

dffeas \phys_cgb[19] (
	.clk(clk),
	.d(ctrl_rdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[19]~q ),
	.prn(vcc));
defparam \phys_cgb[19] .is_wysiwyg = "true";
defparam \phys_cgb[19] .power_up = "low";

dffeas \phys_refclk[19] (
	.clk(clk),
	.d(ctrl_rdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[19]~q ),
	.prn(vcc));
defparam \phys_refclk[19] .is_wysiwyg = "true";
defparam \phys_refclk[19] .power_up = "low";

cyclonev_lcell_comb \modify_data[5]~0 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\mux_pll_type~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\modify_data[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \modify_data[5]~0 .extended_lut = "off";
defparam \modify_data[5]~0 .lut_mask = 64'h2222222222222222;
defparam \modify_data[5]~0 .shared_arith = "off";

dffeas \phys_cgb[0] (
	.clk(clk),
	.d(ctrl_rdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[0]~q ),
	.prn(vcc));
defparam \phys_cgb[0] .is_wysiwyg = "true";
defparam \phys_cgb[0] .power_up = "low";

cyclonev_lcell_comb \uif_rc_sel_wr~0 (
	.dataa(!uif_addr_offset_0),
	.datab(!\uif_cgb_sel_wr~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rc_sel_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rc_sel_wr~0 .extended_lut = "off";
defparam \uif_rc_sel_wr~0 .lut_mask = 64'h2222222222222222;
defparam \uif_rc_sel_wr~0 .shared_arith = "off";

dffeas \pll_uif_rc_sel[2] (
	.clk(clk),
	.d(uif_wdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rc_sel_wr~0_combout ),
	.q(\pll_uif_rc_sel[2]~q ),
	.prn(vcc));
defparam \pll_uif_rc_sel[2] .is_wysiwyg = "true";
defparam \pll_uif_rc_sel[2] .power_up = "low";

cyclonev_lcell_comb \uif_cgb_sel_wr~1 (
	.dataa(!uif_addr_offset_0),
	.datab(!\uif_cgb_sel_wr~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_cgb_sel_wr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_cgb_sel_wr~1 .extended_lut = "off";
defparam \uif_cgb_sel_wr~1 .lut_mask = 64'h1111111111111111;
defparam \uif_cgb_sel_wr~1 .shared_arith = "off";

dffeas \pll_uif_cgb_sel[2] (
	.clk(clk),
	.d(uif_wdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_cgb_sel_wr~1_combout ),
	.q(\pll_uif_cgb_sel[2]~q ),
	.prn(vcc));
defparam \pll_uif_cgb_sel[2] .is_wysiwyg = "true";
defparam \pll_uif_cgb_sel[2] .power_up = "low";

cyclonev_lcell_comb \logical_index[2]~0 (
	.dataa(!\pll_uif_rc_sel[2]~q ),
	.datab(!\pll_uif_cgb_sel[2]~q ),
	.datac(!\mif_req~q ),
	.datad(!\pll_uif_type~q ),
	.datae(!mif_rec_addr_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\logical_index[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \logical_index[2]~0 .extended_lut = "off";
defparam \logical_index[2]~0 .lut_mask = 64'h50305F3F50305F3F;
defparam \logical_index[2]~0 .shared_arith = "off";

dffeas \pll_uif_rc_sel[0] (
	.clk(clk),
	.d(uif_wdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rc_sel_wr~0_combout ),
	.q(\pll_uif_rc_sel[0]~q ),
	.prn(vcc));
defparam \pll_uif_rc_sel[0] .is_wysiwyg = "true";
defparam \pll_uif_rc_sel[0] .power_up = "low";

dffeas \pll_uif_cgb_sel[0] (
	.clk(clk),
	.d(uif_wdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_cgb_sel_wr~1_combout ),
	.q(\pll_uif_cgb_sel[0]~q ),
	.prn(vcc));
defparam \pll_uif_cgb_sel[0] .is_wysiwyg = "true";
defparam \pll_uif_cgb_sel[0] .power_up = "low";

cyclonev_lcell_comb \logical_index[0]~1 (
	.dataa(!\pll_uif_rc_sel[0]~q ),
	.datab(!\pll_uif_cgb_sel[0]~q ),
	.datac(!\mif_req~q ),
	.datad(!\pll_uif_type~q ),
	.datae(!mif_rec_addr_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\logical_index[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \logical_index[0]~1 .extended_lut = "off";
defparam \logical_index[0]~1 .lut_mask = 64'h50305F3F50305F3F;
defparam \logical_index[0]~1 .shared_arith = "off";

dffeas \pll_uif_rc_sel[1] (
	.clk(clk),
	.d(uif_wdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_rc_sel_wr~0_combout ),
	.q(\pll_uif_rc_sel[1]~q ),
	.prn(vcc));
defparam \pll_uif_rc_sel[1] .is_wysiwyg = "true";
defparam \pll_uif_rc_sel[1] .power_up = "low";

dffeas \pll_uif_cgb_sel[1] (
	.clk(clk),
	.d(uif_wdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\uif_cgb_sel_wr~1_combout ),
	.q(\pll_uif_cgb_sel[1]~q ),
	.prn(vcc));
defparam \pll_uif_cgb_sel[1] .is_wysiwyg = "true";
defparam \pll_uif_cgb_sel[1] .power_up = "low";

cyclonev_lcell_comb \logical_index[1]~2 (
	.dataa(!\pll_uif_rc_sel[1]~q ),
	.datab(!\pll_uif_cgb_sel[1]~q ),
	.datac(!\mif_req~q ),
	.datad(!\pll_uif_type~q ),
	.datae(!mif_rec_addr_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\logical_index[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \logical_index[1]~2 .extended_lut = "off";
defparam \logical_index[1]~2 .lut_mask = 64'h50305F3F50305F3F;
defparam \logical_index[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!\logical_index[2]~0_combout ),
	.datab(!\logical_index[0]~1_combout ),
	.datac(!\logical_index[1]~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "off";
defparam \Mux21~0 .lut_mask = 64'h9595959595959595;
defparam \Mux21~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~1 (
	.dataa(!\logical_index[2]~0_combout ),
	.datab(!\logical_index[0]~1_combout ),
	.datac(!\logical_index[1]~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~1 .extended_lut = "off";
defparam \Mux21~1 .lut_mask = 64'h0808080808080808;
defparam \Mux21~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!\phys_cgb[4]~q ),
	.datab(!\phys_cgb[12]~q ),
	.datac(!\phys_cgb[16]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "off";
defparam \Mux23~0 .lut_mask = 64'h000F550000003300;
defparam \Mux23~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux23~1 (
	.dataa(!\phys_cgb[0]~q ),
	.datab(!\phys_cgb[8]~q ),
	.datac(!\Mux21~0_combout ),
	.datad(!\Mux21~1_combout ),
	.datae(!\Mux23~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~1 .extended_lut = "off";
defparam \Mux23~1 .lut_mask = 64'hFACA0000FACA0000;
defparam \Mux23~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!\phys_cgb[7]~q ),
	.datab(!\phys_cgb[15]~q ),
	.datac(!\phys_cgb[19]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "off";
defparam \Mux20~0 .lut_mask = 64'h000F550000003300;
defparam \Mux20~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~1 (
	.dataa(!\phys_cgb[3]~q ),
	.datab(!\phys_cgb[11]~q ),
	.datac(!\logical_index[2]~0_combout ),
	.datad(!\logical_index[0]~1_combout ),
	.datae(!\logical_index[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~1 .extended_lut = "off";
defparam \Mux20~1 .lut_mask = 64'h5005350550053505;
defparam \Mux20~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~2 (
	.dataa(!\Mux20~0_combout ),
	.datab(!\Mux20~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~2 .extended_lut = "off";
defparam \Mux20~2 .lut_mask = 64'h8888888888888888;
defparam \Mux20~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~2 (
	.dataa(!\phys_cgb[6]~q ),
	.datab(!\phys_cgb[14]~q ),
	.datac(!\phys_cgb[18]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~2 .extended_lut = "off";
defparam \Mux21~2 .lut_mask = 64'h000F550000003300;
defparam \Mux21~2 .shared_arith = "off";

dffeas \phys_cgb[2] (
	.clk(clk),
	.d(ctrl_rdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[2]~q ),
	.prn(vcc));
defparam \phys_cgb[2] .is_wysiwyg = "true";
defparam \phys_cgb[2] .power_up = "low";

cyclonev_lcell_comb \Mux21~3 (
	.dataa(!\phys_cgb[2]~q ),
	.datab(!\phys_cgb[10]~q ),
	.datac(!\logical_index[2]~0_combout ),
	.datad(!\logical_index[0]~1_combout ),
	.datae(!\logical_index[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~3 .extended_lut = "off";
defparam \Mux21~3 .lut_mask = 64'h5005350550053505;
defparam \Mux21~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~4 (
	.dataa(!\Mux21~2_combout ),
	.datab(!\Mux21~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~4 .extended_lut = "off";
defparam \Mux21~4 .lut_mask = 64'h8888888888888888;
defparam \Mux21~4 .shared_arith = "off";

cyclonev_lcell_comb \always11~0 (
	.dataa(!ctrl_opcode_2),
	.datab(!ctrl_opcode_0),
	.datac(!waitrequest_to_ctrl),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always11~0 .extended_lut = "off";
defparam \always11~0 .lut_mask = 64'h8080808080808080;
defparam \always11~0 .shared_arith = "off";

dffeas \saved_read_data[1] (
	.clk(clk),
	.d(ctrl_rdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[1]~q ),
	.prn(vcc));
defparam \saved_read_data[1] .is_wysiwyg = "true";
defparam \saved_read_data[1] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~0 (
	.dataa(!\modify_data[5]~0_combout ),
	.datab(!\Mux23~1_combout ),
	.datac(!\Mux20~2_combout ),
	.datad(!\Mux21~4_combout ),
	.datae(!\saved_read_data[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~0 .extended_lut = "off";
defparam \ctrl_wdata~0 .lut_mask = 64'h0004AAAE0004AAAE;
defparam \ctrl_wdata~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata[1]~1 (
	.dataa(!pll_mif_busy1),
	.datab(!\pll_state.PLL_WR~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata[1]~1 .extended_lut = "off";
defparam \ctrl_wdata[1]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ctrl_wdata[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~0 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\pll_state.PLL_RD_L2P~q ),
	.datac(!\mux_pll_type~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~0 .extended_lut = "off";
defparam \ctrl_addr~0 .lut_mask = 64'h4343434343434343;
defparam \ctrl_addr~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~1 (
	.dataa(!\pll_state.PLL_CHK_WORDS~q ),
	.datab(!\pll_state.PLL_DECIDE~q ),
	.datac(!\pll_state.PLL_WAIT~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~1 .extended_lut = "off";
defparam \ctrl_addr~1 .lut_mask = 64'h8080808080808080;
defparam \ctrl_addr~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!\phys_cgb[5]~q ),
	.datab(!\phys_cgb[13]~q ),
	.datac(!\phys_cgb[17]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "off";
defparam \Mux22~0 .lut_mask = 64'h000F550000003300;
defparam \Mux22~0 .shared_arith = "off";

dffeas \phys_cgb[1] (
	.clk(clk),
	.d(ctrl_rdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\phys_cgb[1]~q ),
	.prn(vcc));
defparam \phys_cgb[1] .is_wysiwyg = "true";
defparam \phys_cgb[1] .power_up = "low";

cyclonev_lcell_comb \Mux22~1 (
	.dataa(!\phys_cgb[1]~q ),
	.datab(!\phys_cgb[9]~q ),
	.datac(!\logical_index[2]~0_combout ),
	.datad(!\logical_index[0]~1_combout ),
	.datae(!\logical_index[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~1 .extended_lut = "off";
defparam \Mux22~1 .lut_mask = 64'h5005350550053505;
defparam \Mux22~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux22~2 (
	.dataa(!\Mux22~0_combout ),
	.datab(!\Mux22~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~2 .extended_lut = "off";
defparam \Mux22~2 .lut_mask = 64'h8888888888888888;
defparam \Mux22~2 .shared_arith = "off";

dffeas \saved_read_data[2] (
	.clk(clk),
	.d(ctrl_rdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[2]~q ),
	.prn(vcc));
defparam \saved_read_data[2] .is_wysiwyg = "true";
defparam \saved_read_data[2] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~24 (
	.dataa(!\Mux20~2_combout ),
	.datab(!\Mux21~4_combout ),
	.datac(!\Mux22~2_combout ),
	.datad(!\Mux23~1_combout ),
	.datae(!\saved_read_data[2]~q ),
	.dataf(!\modify_data[5]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~24 .extended_lut = "off";
defparam \ctrl_wdata~24 .lut_mask = 64'h0000FFFFE8ABE8AB;
defparam \ctrl_wdata~24 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~2 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\mux_pll_type~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~2 .extended_lut = "off";
defparam \ctrl_addr~2 .lut_mask = 64'h8888888888888888;
defparam \ctrl_addr~2 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~3 (
	.dataa(!\pll_state.PLL_RD_L2P~q ),
	.datab(!\ctrl_addr~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~3 .extended_lut = "off";
defparam \ctrl_addr~3 .lut_mask = 64'h2222222222222222;
defparam \ctrl_addr~3 .shared_arith = "off";

dffeas \saved_read_data[0] (
	.clk(clk),
	.d(ctrl_rdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[0]~q ),
	.prn(vcc));
defparam \saved_read_data[0] .is_wysiwyg = "true";
defparam \saved_read_data[0] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~2 (
	.dataa(!\saved_read_data[0]~q ),
	.datab(!\modify_data[5]~0_combout ),
	.datac(!\Mux22~2_combout ),
	.datad(!\Mux23~1_combout ),
	.datae(!\Mux20~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~2 .extended_lut = "off";
defparam \ctrl_wdata~2 .lut_mask = 64'h4444474444444744;
defparam \ctrl_wdata~2 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~4 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\pll_state.PLL_RD_L2P~q ),
	.datac(!\mux_pll_type~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~4 .extended_lut = "off";
defparam \ctrl_addr~4 .lut_mask = 64'h3434343434343434;
defparam \ctrl_addr~4 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_addr~5 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\pll_state.PLL_RD_L2P~q ),
	.datac(!\mux_pll_type~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_addr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_addr~5 .extended_lut = "off";
defparam \ctrl_addr~5 .lut_mask = 64'h4040404040404040;
defparam \ctrl_addr~5 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!\Mux23~1_combout ),
	.datab(!\Mux22~2_combout ),
	.datac(!\Mux21~4_combout ),
	.datad(!\Mux20~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'h003A003A003A003A;
defparam \WideOr1~0 .shared_arith = "off";

dffeas \saved_read_data[5] (
	.clk(clk),
	.d(ctrl_rdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[5]~q ),
	.prn(vcc));
defparam \saved_read_data[5] .is_wysiwyg = "true";
defparam \saved_read_data[5] .power_up = "low";

dffeas \phys_refclk[2] (
	.clk(clk),
	.d(ctrl_rdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[2]~q ),
	.prn(vcc));
defparam \phys_refclk[2] .is_wysiwyg = "true";
defparam \phys_refclk[2] .power_up = "low";

dffeas \phys_refclk[22] (
	.clk(clk),
	.d(readdata_for_user_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[22]~q ),
	.prn(vcc));
defparam \phys_refclk[22] .is_wysiwyg = "true";
defparam \phys_refclk[22] .power_up = "low";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!\phys_refclk[7]~q ),
	.datab(!\phys_refclk[17]~q ),
	.datac(!\phys_refclk[22]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "off";
defparam \Mux26~0 .lut_mask = 64'h000F550000003300;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~1 (
	.dataa(!\phys_refclk[2]~q ),
	.datab(!\phys_refclk[12]~q ),
	.datac(!\Mux21~0_combout ),
	.datad(!\Mux21~1_combout ),
	.datae(!\Mux26~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~1 .extended_lut = "off";
defparam \Mux26~1 .lut_mask = 64'h0535FFFF0535FFFF;
defparam \Mux26~1 .shared_arith = "off";

dffeas \phys_refclk[23] (
	.clk(clk),
	.d(readdata_for_user_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[23]~q ),
	.prn(vcc));
defparam \phys_refclk[23] .is_wysiwyg = "true";
defparam \phys_refclk[23] .power_up = "low";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!\phys_refclk[8]~q ),
	.datab(!\phys_refclk[18]~q ),
	.datac(!\phys_refclk[23]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "off";
defparam \Mux25~0 .lut_mask = 64'h000F550000003300;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~1 (
	.dataa(!\phys_refclk[3]~q ),
	.datab(!\phys_refclk[13]~q ),
	.datac(!\Mux21~0_combout ),
	.datad(!\Mux21~1_combout ),
	.datae(!\Mux25~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~1 .extended_lut = "off";
defparam \Mux25~1 .lut_mask = 64'h0535FFFF0535FFFF;
defparam \Mux25~1 .shared_arith = "off";

dffeas \phys_refclk[1] (
	.clk(clk),
	.d(ctrl_rdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[1]~q ),
	.prn(vcc));
defparam \phys_refclk[1] .is_wysiwyg = "true";
defparam \phys_refclk[1] .power_up = "low";

dffeas \phys_refclk[21] (
	.clk(clk),
	.d(readdata_for_user_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[21]~q ),
	.prn(vcc));
defparam \phys_refclk[21] .is_wysiwyg = "true";
defparam \phys_refclk[21] .power_up = "low";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!\phys_refclk[6]~q ),
	.datab(!\phys_refclk[16]~q ),
	.datac(!\phys_refclk[21]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "off";
defparam \Mux27~0 .lut_mask = 64'h000F550000003300;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~1 (
	.dataa(!\phys_refclk[1]~q ),
	.datab(!\phys_refclk[11]~q ),
	.datac(!\Mux21~0_combout ),
	.datad(!\Mux21~1_combout ),
	.datae(!\Mux27~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~1 .extended_lut = "off";
defparam \Mux27~1 .lut_mask = 64'h0535FFFF0535FFFF;
defparam \Mux27~1 .shared_arith = "off";

dffeas \phys_refclk[0] (
	.clk(clk),
	.d(ctrl_rdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[0]~q ),
	.prn(vcc));
defparam \phys_refclk[0] .is_wysiwyg = "true";
defparam \phys_refclk[0] .power_up = "low";

dffeas \phys_refclk[20] (
	.clk(clk),
	.d(readdata_for_user_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[20]~q ),
	.prn(vcc));
defparam \phys_refclk[20] .is_wysiwyg = "true";
defparam \phys_refclk[20] .power_up = "low";

cyclonev_lcell_comb \Mux28~0 (
	.dataa(!\phys_refclk[5]~q ),
	.datab(!\phys_refclk[15]~q ),
	.datac(!\phys_refclk[20]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~0 .extended_lut = "off";
defparam \Mux28~0 .lut_mask = 64'h000F550000003300;
defparam \Mux28~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~1 (
	.dataa(!\phys_refclk[0]~q ),
	.datab(!\phys_refclk[10]~q ),
	.datac(!\Mux21~0_combout ),
	.datad(!\Mux21~1_combout ),
	.datae(!\Mux28~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~1 .extended_lut = "off";
defparam \Mux28~1 .lut_mask = 64'h0535FFFF0535FFFF;
defparam \Mux28~1 .shared_arith = "off";

dffeas \phys_refclk[24] (
	.clk(clk),
	.d(readdata_for_user_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\phys_refclk[0]~0_combout ),
	.q(\phys_refclk[24]~q ),
	.prn(vcc));
defparam \phys_refclk[24] .is_wysiwyg = "true";
defparam \phys_refclk[24] .power_up = "low";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!\phys_refclk[9]~q ),
	.datab(!\phys_refclk[19]~q ),
	.datac(!\phys_refclk[24]~q ),
	.datad(!\logical_index[2]~0_combout ),
	.datae(!\logical_index[0]~1_combout ),
	.dataf(!\logical_index[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "off";
defparam \Mux24~0 .lut_mask = 64'h000F550000003300;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~1 (
	.dataa(!\phys_refclk[4]~q ),
	.datab(!\phys_refclk[14]~q ),
	.datac(!\Mux21~0_combout ),
	.datad(!\Mux21~1_combout ),
	.datae(!\Mux24~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~1 .extended_lut = "off";
defparam \Mux24~1 .lut_mask = 64'h0535FFFF0535FFFF;
defparam \Mux24~1 .shared_arith = "off";

cyclonev_lcell_comb \modify_data[5]~1 (
	.dataa(!\Mux26~1_combout ),
	.datab(!\Mux25~1_combout ),
	.datac(!\Mux27~1_combout ),
	.datad(!\Mux28~1_combout ),
	.datae(!\Mux24~1_combout ),
	.dataf(!\ctrl_addr~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\modify_data[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \modify_data[5]~1 .extended_lut = "off";
defparam \modify_data[5]~1 .lut_mask = 64'h0000000044482000;
defparam \modify_data[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \modify_data[5]~2 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\mux_pll_type~0_combout ),
	.datac(!\WideOr1~0_combout ),
	.datad(!\saved_read_data[5]~q ),
	.datae(!\modify_data[5]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\modify_data[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \modify_data[5]~2 .extended_lut = "off";
defparam \modify_data[5]~2 .lut_mask = 64'h2031FFFF2031FFFF;
defparam \modify_data[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \Ram0~3 (
	.dataa(!\Mux27~1_combout ),
	.datab(!\Mux26~1_combout ),
	.datac(!\Mux25~1_combout ),
	.datad(!\Mux24~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Ram0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Ram0~3 .extended_lut = "off";
defparam \Ram0~3 .lut_mask = 64'h0180018001800180;
defparam \Ram0~3 .shared_arith = "off";

dffeas \saved_read_data[3] (
	.clk(clk),
	.d(ctrl_rdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[3]~q ),
	.prn(vcc));
defparam \saved_read_data[3] .is_wysiwyg = "true";
defparam \saved_read_data[3] .power_up = "low";

dffeas \saved_read_data[9] (
	.clk(clk),
	.d(ctrl_rdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[9]~q ),
	.prn(vcc));
defparam \saved_read_data[9] .is_wysiwyg = "true";
defparam \saved_read_data[9] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!\Mux22~0_combout ),
	.datab(!\Mux20~0_combout ),
	.datac(!\Mux22~1_combout ),
	.datad(!\Mux20~1_combout ),
	.datae(!\Mux21~2_combout ),
	.dataf(!\Mux21~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h20A04C004C004C00;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \modify_data[9]~3 (
	.dataa(!\Ram0~3_combout ),
	.datab(!\saved_read_data[3]~q ),
	.datac(!\saved_read_data[9]~q ),
	.datad(!\WideOr0~0_combout ),
	.datae(!\word_cnt[0]~q ),
	.dataf(!\mux_pll_type~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\modify_data[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \modify_data[9]~3 .extended_lut = "off";
defparam \modify_data[9]~3 .lut_mask = 64'h555533330F0F00FF;
defparam \modify_data[9]~3 .shared_arith = "off";

dffeas \saved_read_data[13] (
	.clk(clk),
	.d(ctrl_rdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[13]~q ),
	.prn(vcc));
defparam \saved_read_data[13] .is_wysiwyg = "true";
defparam \saved_read_data[13] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~17 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\mux_pll_type~0_combout ),
	.datac(!\saved_read_data[1]~q ),
	.datad(!\saved_read_data[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~17 .extended_lut = "off";
defparam \ctrl_wdata~17 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \ctrl_wdata~17 .shared_arith = "off";

dffeas \saved_read_data[14] (
	.clk(clk),
	.d(ctrl_rdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[14]~q ),
	.prn(vcc));
defparam \saved_read_data[14] .is_wysiwyg = "true";
defparam \saved_read_data[14] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~18 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\mux_pll_type~0_combout ),
	.datac(!\saved_read_data[2]~q ),
	.datad(!\saved_read_data[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~18 .extended_lut = "off";
defparam \ctrl_wdata~18 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \ctrl_wdata~18 .shared_arith = "off";

dffeas \saved_read_data[15] (
	.clk(clk),
	.d(ctrl_rdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[15]~q ),
	.prn(vcc));
defparam \saved_read_data[15] .is_wysiwyg = "true";
defparam \saved_read_data[15] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~19 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\mux_pll_type~0_combout ),
	.datac(!\saved_read_data[3]~q ),
	.datad(!\saved_read_data[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~19 .extended_lut = "off";
defparam \ctrl_wdata~19 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \ctrl_wdata~19 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~2 (
	.dataa(!\word_cnt[0]~q ),
	.datab(!\pll_state.PLL_CHK_WORDS~q ),
	.datac(!\uif_l2p_active~q ),
	.datad(!waitrequest_to_ctrl),
	.datae(!\pll_state.PLL_DECIDE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~2 .extended_lut = "off";
defparam \Selector0~2 .lut_mask = 64'h22222F2222222F22;
defparam \Selector0~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~3 (
	.dataa(!pll_mif_busy1),
	.datab(!pll_go),
	.datac(!\pll_uif_go~q ),
	.datad(!\always13~0_combout ),
	.datae(!\Selector0~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~3 .extended_lut = "off";
defparam \Selector0~3 .lut_mask = 64'h7FFF00007FFF0000;
defparam \Selector0~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!\pll_uif_cgb_sel[0]~q ),
	.datab(!\phys_cgb[0]~q ),
	.datac(!\phys_refclk[0]~q ),
	.datad(!uif_addr_offset_0),
	.datae(!uif_addr_offset_1),
	.dataf(!uif_addr_offset_2),
	.datag(!\pll_uif_rc_sel[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "on";
defparam \Mux19~0 .lut_mask = 64'h0F550F3300000000;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!\pll_uif_cgb_sel[1]~q ),
	.datab(!\phys_cgb[1]~q ),
	.datac(!\phys_refclk[1]~q ),
	.datad(!uif_addr_offset_0),
	.datae(!uif_addr_offset_1),
	.dataf(!uif_addr_offset_2),
	.datag(!\pll_uif_rc_sel[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "on";
defparam \Mux18~0 .lut_mask = 64'h0F550F3300000000;
defparam \Mux18~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!\pll_uif_cgb_sel[2]~q ),
	.datab(!\phys_cgb[2]~q ),
	.datac(!\phys_refclk[2]~q ),
	.datad(!uif_addr_offset_0),
	.datae(!uif_addr_offset_1),
	.dataf(!uif_addr_offset_2),
	.datag(!\pll_uif_rc_sel[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "on";
defparam \Mux17~0 .lut_mask = 64'h0F550F3300000000;
defparam \Mux17~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~0 (
	.dataa(!uif_addr_offset_0),
	.datab(!\Equal3~0_combout ),
	.datac(!\phys_refclk[20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~0 .extended_lut = "off";
defparam \uif_rdata~0 .lut_mask = 64'h0808080808080808;
defparam \uif_rdata~0 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~1 (
	.dataa(!uif_addr_offset_0),
	.datab(!\Equal3~0_combout ),
	.datac(!\phys_refclk[21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~1 .extended_lut = "off";
defparam \uif_rdata~1 .lut_mask = 64'h0808080808080808;
defparam \uif_rdata~1 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~2 (
	.dataa(!uif_addr_offset_0),
	.datab(!\Equal3~0_combout ),
	.datac(!\phys_refclk[22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~2 .extended_lut = "off";
defparam \uif_rdata~2 .lut_mask = 64'h0808080808080808;
defparam \uif_rdata~2 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~3 (
	.dataa(!uif_addr_offset_0),
	.datab(!\Equal3~0_combout ),
	.datac(!\phys_refclk[23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~3 .extended_lut = "off";
defparam \uif_rdata~3 .lut_mask = 64'h0808080808080808;
defparam \uif_rdata~3 .shared_arith = "off";

cyclonev_lcell_comb \uif_rdata~4 (
	.dataa(!uif_addr_offset_0),
	.datab(!\Equal3~0_combout ),
	.datac(!\phys_refclk[24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\uif_rdata~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \uif_rdata~4 .extended_lut = "off";
defparam \uif_rdata~4 .lut_mask = 64'h0808080808080808;
defparam \uif_rdata~4 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_lock~0 (
	.dataa(!pll_mif_busy1),
	.datab(!\uif_l2p_active~q ),
	.datac(!\state_event[1]~q ),
	.datad(!\state_event[0]~q ),
	.datae(!\state_event[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_lock~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_lock~0 .extended_lut = "off";
defparam \ctrl_lock~0 .lut_mask = 64'h4440000044400000;
defparam \ctrl_lock~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode[0]~0 (
	.dataa(!\ctrl_go~0_combout ),
	.datab(!\Selector0~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode[0]~0 .extended_lut = "off";
defparam \ctrl_opcode[0]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \ctrl_opcode[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_opcode~1 (
	.dataa(!\pll_state.PLL_RD_L2P~q ),
	.datab(!\pll_state.PLL_RD~q ),
	.datac(!\Selector0~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_opcode~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_opcode~1 .extended_lut = "off";
defparam \ctrl_opcode~1 .lut_mask = 64'h0808080808080808;
defparam \ctrl_opcode~1 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~3 (
	.dataa(!\Mux26~1_combout ),
	.datab(!\Mux25~1_combout ),
	.datac(!\Mux27~1_combout ),
	.datad(!\Mux28~1_combout ),
	.datae(!\Mux24~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~3 .extended_lut = "off";
defparam \ctrl_wdata~3 .lut_mask = 64'hEE001313EE001313;
defparam \ctrl_wdata~3 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata[4]~4 (
	.dataa(!pll_mif_busy1),
	.datab(!\ctrl_addr~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata[4]~4 .extended_lut = "off";
defparam \ctrl_wdata[4]~4 .lut_mask = 64'h4444444444444444;
defparam \ctrl_wdata[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata[4]~5 (
	.dataa(!pll_mif_busy1),
	.datab(!\modify_data[5]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata[4]~5 .extended_lut = "off";
defparam \ctrl_wdata[4]~5 .lut_mask = 64'h4444444444444444;
defparam \ctrl_wdata[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \WideOr2~0 (
	.dataa(!\Mux23~1_combout ),
	.datab(!\Mux22~2_combout ),
	.datac(!\Mux21~4_combout ),
	.datad(!\Mux20~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr2~0 .extended_lut = "off";
defparam \WideOr2~0 .lut_mask = 64'h01BE01BE01BE01BE;
defparam \WideOr2~0 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~6 (
	.dataa(!\ctrl_wdata~3_combout ),
	.datab(!\ctrl_wdata[4]~4_combout ),
	.datac(!\ctrl_wdata[4]~5_combout ),
	.datad(!\saved_read_data[3]~q ),
	.datae(!\WideOr2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~6 .extended_lut = "off";
defparam \ctrl_wdata~6 .lut_mask = 64'h3437040734370407;
defparam \ctrl_wdata~6 .shared_arith = "off";

cyclonev_lcell_comb \Ram0~0 (
	.dataa(!\Mux28~1_combout ),
	.datab(!\Mux27~1_combout ),
	.datac(!\Mux26~1_combout ),
	.datad(!\Mux25~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Ram0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Ram0~0 .extended_lut = "off";
defparam \Ram0~0 .lut_mask = 64'h6660666066606660;
defparam \Ram0~0 .shared_arith = "off";

dffeas \saved_read_data[4] (
	.clk(clk),
	.d(ctrl_rdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[4]~q ),
	.prn(vcc));
defparam \saved_read_data[4] .is_wysiwyg = "true";
defparam \saved_read_data[4] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~7 (
	.dataa(!\Mux24~1_combout ),
	.datab(!\ctrl_wdata[4]~4_combout ),
	.datac(!\ctrl_wdata[4]~5_combout ),
	.datad(!\Ram0~0_combout ),
	.datae(!\saved_read_data[4]~q ),
	.dataf(!\WideOr1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~7 .extended_lut = "off";
defparam \ctrl_wdata~7 .lut_mask = 64'h0008030B3038333B;
defparam \ctrl_wdata~7 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~8 (
	.dataa(!\Mux26~1_combout ),
	.datab(!\Mux25~1_combout ),
	.datac(!\Mux27~1_combout ),
	.datad(!\Mux28~1_combout ),
	.datae(!\Mux24~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~8 .extended_lut = "off";
defparam \ctrl_wdata~8 .lut_mask = 64'h2224200022242000;
defparam \ctrl_wdata~8 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata[6]~9 (
	.dataa(!pll_mif_busy1),
	.datab(!\word_cnt[0]~q ),
	.datac(!\mux_pll_type~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata[6]~9 .extended_lut = "off";
defparam \ctrl_wdata[6]~9 .lut_mask = 64'hBABABABABABABABA;
defparam \ctrl_wdata[6]~9 .shared_arith = "off";

dffeas \saved_read_data[6] (
	.clk(clk),
	.d(ctrl_rdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[6]~q ),
	.prn(vcc));
defparam \saved_read_data[6] .is_wysiwyg = "true";
defparam \saved_read_data[6] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~10 (
	.dataa(!\saved_read_data[0]~q ),
	.datab(!\ctrl_wdata[4]~4_combout ),
	.datac(!\ctrl_wdata~8_combout ),
	.datad(!\ctrl_wdata[6]~9_combout ),
	.datae(!\saved_read_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~10 .extended_lut = "off";
defparam \ctrl_wdata~10 .lut_mask = 64'h0C113F110C113F11;
defparam \ctrl_wdata~10 .shared_arith = "off";

cyclonev_lcell_comb \Ram0~1 (
	.dataa(!\Mux24~1_combout ),
	.datab(!\Mux27~1_combout ),
	.datac(!\Mux26~1_combout ),
	.datad(!\Mux25~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Ram0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Ram0~1 .extended_lut = "off";
defparam \Ram0~1 .lut_mask = 64'h542A542A542A542A;
defparam \Ram0~1 .shared_arith = "off";

dffeas \saved_read_data[7] (
	.clk(clk),
	.d(ctrl_rdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[7]~q ),
	.prn(vcc));
defparam \saved_read_data[7] .is_wysiwyg = "true";
defparam \saved_read_data[7] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~11 (
	.dataa(!\Mux28~1_combout ),
	.datab(!\ctrl_wdata[4]~4_combout ),
	.datac(!\saved_read_data[1]~q ),
	.datad(!\ctrl_wdata[6]~9_combout ),
	.datae(!\Ram0~1_combout ),
	.dataf(!\saved_read_data[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~11 .extended_lut = "off";
defparam \ctrl_wdata~11 .lut_mask = 64'h0003440333037703;
defparam \ctrl_wdata~11 .shared_arith = "off";

cyclonev_lcell_comb \Ram0~2 (
	.dataa(!\Mux27~1_combout ),
	.datab(!\Mux26~1_combout ),
	.datac(!\Mux25~1_combout ),
	.datad(!\Mux24~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Ram0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Ram0~2 .extended_lut = "off";
defparam \Ram0~2 .lut_mask = 64'h02A002A002A002A0;
defparam \Ram0~2 .shared_arith = "off";

dffeas \saved_read_data[8] (
	.clk(clk),
	.d(ctrl_rdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[8]~q ),
	.prn(vcc));
defparam \saved_read_data[8] .is_wysiwyg = "true";
defparam \saved_read_data[8] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~12 (
	.dataa(!\ctrl_wdata[4]~4_combout ),
	.datab(!\saved_read_data[2]~q ),
	.datac(!\ctrl_wdata[6]~9_combout ),
	.datad(!\Ram0~2_combout ),
	.datae(!\saved_read_data[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~12 .extended_lut = "off";
defparam \ctrl_wdata~12 .lut_mask = 64'h01A151F101A151F1;
defparam \ctrl_wdata~12 .shared_arith = "off";

cyclonev_lcell_comb \Ram0~4 (
	.dataa(!\Mux27~1_combout ),
	.datab(!\Mux26~1_combout ),
	.datac(!\Mux25~1_combout ),
	.datad(!\Mux24~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Ram0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Ram0~4 .extended_lut = "off";
defparam \Ram0~4 .lut_mask = 64'h0060006000600060;
defparam \Ram0~4 .shared_arith = "off";

dffeas \saved_read_data[10] (
	.clk(clk),
	.d(ctrl_rdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[10]~q ),
	.prn(vcc));
defparam \saved_read_data[10] .is_wysiwyg = "true";
defparam \saved_read_data[10] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~13 (
	.dataa(!\ctrl_wdata[4]~4_combout ),
	.datab(!\saved_read_data[4]~q ),
	.datac(!\ctrl_wdata[6]~9_combout ),
	.datad(!\Ram0~4_combout ),
	.datae(!\saved_read_data[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~13 .extended_lut = "off";
defparam \ctrl_wdata~13 .lut_mask = 64'h01A151F101A151F1;
defparam \ctrl_wdata~13 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~14 (
	.dataa(!\Mux22~2_combout ),
	.datab(!\Mux20~2_combout ),
	.datac(!\ctrl_wdata[4]~5_combout ),
	.datad(!\Mux21~4_combout ),
	.datae(!\ctrl_wdata[6]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~14 .extended_lut = "off";
defparam \ctrl_wdata~14 .lut_mask = 64'h2000000020000000;
defparam \ctrl_wdata~14 .shared_arith = "off";

dffeas \saved_read_data[11] (
	.clk(clk),
	.d(ctrl_rdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[11]~q ),
	.prn(vcc));
defparam \saved_read_data[11] .is_wysiwyg = "true";
defparam \saved_read_data[11] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~20 (
	.dataa(!\Mux27~1_combout ),
	.datab(!\Mux25~1_combout ),
	.datac(!\Mux24~1_combout ),
	.datad(!\Mux26~1_combout ),
	.datae(!\ctrl_wdata[6]~9_combout ),
	.dataf(!\Mux28~1_combout ),
	.datag(!\saved_read_data[11]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~20 .extended_lut = "on";
defparam \ctrl_wdata~20 .lut_mask = 64'h0F0F00040F0F0000;
defparam \ctrl_wdata~20 .shared_arith = "off";

cyclonev_lcell_comb \ctrl_wdata~15 (
	.dataa(!\Mux23~1_combout ),
	.datab(!\ctrl_wdata[4]~5_combout ),
	.datac(!\ctrl_wdata~14_combout ),
	.datad(!\ctrl_wdata~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~15 .extended_lut = "off";
defparam \ctrl_wdata~15 .lut_mask = 64'h0A3B0A3B0A3B0A3B;
defparam \ctrl_wdata~15 .shared_arith = "off";

dffeas \saved_read_data[12] (
	.clk(clk),
	.d(ctrl_rdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\saved_read_data[12]~q ),
	.prn(vcc));
defparam \saved_read_data[12] .is_wysiwyg = "true";
defparam \saved_read_data[12] .power_up = "low";

cyclonev_lcell_comb \ctrl_wdata~16 (
	.dataa(!\saved_read_data[0]~q ),
	.datab(!\Mux23~1_combout ),
	.datac(!\ctrl_wdata[4]~5_combout ),
	.datad(!\ctrl_wdata[6]~9_combout ),
	.datae(!\ctrl_wdata~14_combout ),
	.dataf(!\saved_read_data[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctrl_wdata~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_wdata~16 .extended_lut = "off";
defparam \ctrl_wdata~16 .lut_mask = 64'h000533370F053F37;
defparam \ctrl_wdata~16 .shared_arith = "off";

endmodule

module RECONFIGURE_IP_alt_xcvr_resync_4 (
	resync_chains0sync_r_1,
	clk,
	mgmt_rst_reset)/* synthesis synthesis_greybox=0 */;
output 	resync_chains0sync_r_1;
input 	clk;
input 	mgmt_rst_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \resync_chains[0].sync_r[0]~0_combout ;
wire \resync_chains[0].sync_r[0]~q ;


dffeas \resync_chains[0].sync_r[1] (
	.clk(clk),
	.d(\resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resync_chains0sync_r_1),
	.prn(vcc));
defparam \resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[1] .power_up = "low";

cyclonev_lcell_comb \resync_chains[0].sync_r[0]~0 (
	.dataa(!mgmt_rst_reset),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\resync_chains[0].sync_r[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \resync_chains[0].sync_r[0]~0 .extended_lut = "off";
defparam \resync_chains[0].sync_r[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \resync_chains[0].sync_r[0]~0 .shared_arith = "off";

dffeas \resync_chains[0].sync_r[0] (
	.clk(clk),
	.d(\resync_chains[0].sync_r[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[0] .power_up = "low";

endmodule
