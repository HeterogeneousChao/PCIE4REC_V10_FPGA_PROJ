// RECONFIGURE_IP.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module RECONFIGURE_IP (
		output wire        reconfig_busy,             //      reconfig_busy.reconfig_busy
		input  wire        mgmt_clk_clk,              //       mgmt_clk_clk.clk
		input  wire        mgmt_rst_reset,            //     mgmt_rst_reset.reset
		input  wire [6:0]  reconfig_mgmt_address,     //      reconfig_mgmt.address
		input  wire        reconfig_mgmt_read,        //                   .read
		output wire [31:0] reconfig_mgmt_readdata,    //                   .readdata
		output wire        reconfig_mgmt_waitrequest, //                   .waitrequest
		input  wire        reconfig_mgmt_write,       //                   .write
		input  wire [31:0] reconfig_mgmt_writedata,   //                   .writedata
		output wire [31:0] reconfig_mif_address,      //       reconfig_mif.address
		output wire        reconfig_mif_read,         //                   .read
		input  wire [15:0] reconfig_mif_readdata,     //                   .readdata
		input  wire        reconfig_mif_waitrequest,  //                   .waitrequest
		output wire [69:0] reconfig_to_xcvr,          //   reconfig_to_xcvr.reconfig_to_xcvr
		input  wire [45:0] reconfig_from_xcvr         // reconfig_from_xcvr.reconfig_from_xcvr
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Cyclone V"),
		.number_of_reconfig_interfaces (1),
		.enable_offset                 (1),
		.enable_lc                     (0),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (1),
		.enable_pll                    (1)
	) reconfigure_ip_inst (
		.reconfig_busy             (reconfig_busy),             //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (mgmt_clk_clk),              //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (mgmt_rst_reset),            //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (reconfig_mgmt_address),     //      reconfig_mgmt.address
		.reconfig_mgmt_read        (reconfig_mgmt_read),        //                   .read
		.reconfig_mgmt_readdata    (reconfig_mgmt_readdata),    //                   .readdata
		.reconfig_mgmt_waitrequest (reconfig_mgmt_waitrequest), //                   .waitrequest
		.reconfig_mgmt_write       (reconfig_mgmt_write),       //                   .write
		.reconfig_mgmt_writedata   (reconfig_mgmt_writedata),   //                   .writedata
		.reconfig_mif_address      (reconfig_mif_address),      //       reconfig_mif.address
		.reconfig_mif_read         (reconfig_mif_read),         //                   .read
		.reconfig_mif_readdata     (reconfig_mif_readdata),     //                   .readdata
		.reconfig_mif_waitrequest  (reconfig_mif_waitrequest),  //                   .waitrequest
		.reconfig_to_xcvr          (reconfig_to_xcvr),          //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (reconfig_from_xcvr),        // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                          //        (terminated)
		.rx_cal_busy               (),                          //        (terminated)
		.cal_busy_in               (1'b0)                       //        (terminated)
	);

endmodule
