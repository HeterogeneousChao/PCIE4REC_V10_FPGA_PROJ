// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:17 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rk8su2FIqu8CSS+3sQzDcmHjt2+Jyf0rr+gjwRVQZwtRDpKz5PHhCiKK8AtFacpH
abw570ju0s2RhwgvMgt4C07hupdbaBo/iqF06tw2zb5px3z5/HNMF5v7Mxy5o/zW
g1WjRqqX7archUSZ8aJQixbPisEqe4unSR8DTR1MzQ4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6544)
FBR1Uz5Ss/yOP/kwXNtfXizmiKDKrpTJG6PMhtri6u37G8GinlBL/s0gAx1YRDID
NSX2x+oj8SKZFExblYutTIU9KQvTnHuDABe+fxxvduC7K7wDaDdwGtNIO5TBQAxu
vycwecNdUs6pjTOLgLJuKSmxIJblkkm171cEkX3HiqQtBb9DRUdACpZmWd1V48CE
e1xQvAsK9CG9zlvUePepE4tVTA8agPdlZK+vTOu5VYOWKMILXdprffO/jf0FvuVP
RsX8awcW9HBYW4YGWl6r2taOOD6j6OChNGAJl/3S3UT4ktlos9kB7XwyEpP6mfFc
nMKZVduFHeIisfogXiH5tD/1iFZQcii1AIrrYtFDIVPaMjc8SQdOXSqba6BGoOLH
C9Cgl4o15miHzuoNJXMdMT/ofTH2iT6NzK4LJf1v5OK4wcGXk/ebHE/QCwc0UJSQ
BYBmqL82DAu2JKYxBw2xROfCqSpI51gH+MUWuzthYNfteowwff4NYeV32//qEN+R
sIYst2tq+1OgqMhUzHHv3Cxti7hubfjk0dbjvUKvuCGTVElvUsLllWKCtTV/hjPp
zspRhb7J2Fr/xZDzaBPa+5HLu9ivGlKkQIyPRQ1nO5V2y6dp51Dvt6EQObK3S0tI
/1wIZoJW9We0CBbk8xbBXFHnTxh5SdHxTizkwP/GfJejyW5t0MM7AoVdvUAWEx0S
tqhPVMQ6cWN6/CiDo8PV0xJHoYVhW2LukfKVQisY7nuGRByJBwSJ37msTk+Z567f
S6xISfXbwj2whV2SpG8mGhmE2WHkdKi1pKqGyuBiBWcdzKYfL7x0ca4cU4PXFnpz
CeJDnDug0kubvN9TBx+fzo6BpzY3k58itXiYPIGZfw3HMmvDzpT+FVbo7EIq5RMX
QjQocMFsGlrcCuaaGrPmGdV5hFrCInoP1o/Du12tsp2X2TACf74o63UrXiISMz91
+Sm0iw+UPME4yu8TgTXXh31h17IBDw/HIbVsVifFPbJw2P0YezaKLEKq1yXhy/Jj
ia/VWVYCMlBZLdYoGJ4S8TPvby32n/CWUA7hH8dayM6M2sPR0UlAEfKRiT82P63W
iZJakd2d2ewksKAi5z4zrjTjPolhVFJDDxwXdr5Y8YVpmE+bP/viJNZVGXYeeBQB
8+8jmOYbKh0lodt1AhR0yAp5DrOdiUHw5FATvvJ51v5npqGUTXQkSX3iBqY8zA++
Q4LbjHgE1YBE1ffIKKCJPUzpS6Eemx2KynMN0CIKkqdB0dDyDBxu4Zv/JBuaNySc
+YPLYiA51oiwYNYb22YB4rUdPtL45CRBfkCSq56kwlH/eBJobBpP/6D44TzuzgMX
fz0DyFs3ifDNH03TyP5/M1tuHFEmZF0Zn5MlQjlEstCzFp5dvVksGAbmqnY0bKsc
PCkw2LZka3UQHIMJzgv+VPZQr9FYvzGEMP6Cib/Eln3i8uI6mYJbEBfDU4Uy+AOc
2uITx4hjYwiPf9RHUmBYIBt0WTEg8Qb/r97IIiAd2oGSv4nqLdI88gE89Vvx1Hil
AB4/xyHambXiVEEkNMG1DxQLacZzS6mOEMx1Uo9a0XAAe4GtdfnwxMhLcqPZqRqi
7MnBdChgw3Ez16mbM98kPLDxfQX2XVcxgR9V6pCRu1C5k1XdDC4fWA78ddJwtpKF
2DDpRfQdWNPT1jky6hx7T+A2sP/3Q/4Cxo9SsdozigIu0bUkxR8XwqkOgLV8p4Qc
dwK4XuALBTjNROexCCMcng+G5NgBgFLtZIDc26kwK/aGVoGHpo4J0P9+Vd3RwgAs
LGpBsyyXsfNwAE4Q0Z+rWzmKxZRlk8XqNdjKgEOFd1IY3zRVvkWjJDuud8FhO5ql
DbxJvqsFa+mlCK4tOqSuVNeVnWKQ4uraek0tpJK8od6xP8uqM1zJ3SPD3mhmlOoa
NTvOUU9COtMedgU5coSNnjKQx8PyZiga5qVX2lk1HA5ISKanPQEcFMZo9hkxKyvl
WOlDDP5+XtIfzmmzGR36tvh8115Fuam6AWdI2KPecKizXMQhJMSpegbRI2Em5kT2
PidpXDWbWBLmQkHX+jNVSp3XXPtqjeRLGzNf3f4pu3wOOoNX/UjY7Yr5/wgtDmYE
yK/NHcAxXS1gniOfPmf6DHSgpeOsn1Q9pSZKM29M7em9QiS0hP33oPsh/eGwJu9X
g7pv80dt8tK4L8Z9g8xZatI50MwXZ/Joyc/oT4U0ovtDKiwgZYpjzJ+DWXbN8Tgx
/iJMOHy2OSKjPtO3BopWPmTXNFCjU0x22ArDNeetlm7c3Mp7GeL+zoGn1uIIEuyt
Y32Ni84jnvdxg/3FKiasxtWqboOSxzoS2paMAoQSzM1pUafu8vvz9tz72SLdlw8P
lc6JjUui1gdsHeSSg5GtBTrHU16fr6DwlsyPI8erSG1csaR3Z/3kAmkydWkF7Uyy
aI1tDZBigbdONFlkTyNE0MejhlqtDl6aDW/zQAa3915ARe9+xHZfw6qGo7Wvddwk
kMTrlaDPHC6F1pzGVjQsZC7JxsZXZQy7BTfe+y9BX80WDNt1IBsL+OT3rTW4w7Mw
92axWkqkwGNXcqV5yXICMslYxgDDB+pYCLCBAxk/WPXjwcOjgWi0+qbqJBCM+B6W
ZiyBAkCrDDQyVFNqikW3CEv30/aJzGJKsFANCci12h9DtakVEKLA3todxHuh+Dj/
zOtWyhhcOchyhhR7B9uY5aiZXvt6IHFBYSeX5ORNkVXC5Ypj7Uh+CFeF3pOwruEl
MTB/BhgUoAMe+X2Gb5IF4dfbDh2d4kn74D2BXK6+dH0PZ5UJ6lituiV23wYS2TQT
h2W1K5Xu1wEM4hiKcSrqu/5PT+QvBMmRPEP+5itNCH0jiPCeknLlZohLdw3WKnhb
+oglfJxPWSMRVrtmeSYdPSKaKKHyXiPQCAc9iccSb5WDyJpxKGKPfA+B43Vzm8Si
c9wWr+m76RygDG+7/gZwDnsC3IXWgBdG5AS1uKI7SEv3W7BMrSOLoeYFJi+lVtmq
rv158q3UdNv2V0ZYUU5ULkqnQo3Obt1JK+as7hHNaQY88WwgDSbp/ej2Ggj94rdm
uCKJFLXHe4ac1pzgdqSSPc+9yV+AQx9uoopqHYkhPU9R1aameCwCexL9BJmdmGml
jbLi6mQKNB//kmyLqMj3cGmDWxY/eqkTzw31AG1NcTLAijbUavak8jAhVWIwlsBS
TZ8xqN3N6Ov+frHrRCUP/76jq9KOFd8WHyMHuDGkWp/GpYjXxujx74WTkyjxsO8v
YP3PLxHXAccvtktsmpIzQv72vFANYDapwKr5pHSRdaD9woLqWmIJwbmBuipH7VaY
aZ0QU3Idc6EHUb9TlvGtGvSXF51TlL6X30dbFls4p42tg5N87DQUqN2KrsQj8bfP
d7rgg1xB0nYWHe1NTzt8qoGn21gS6uUIfdvEncG5vPukHmWxIV1Og4TObTFQ9+zY
Fbof31Xa+7u7oX2UTthjfCzehpi9uFSwjjyIYOHulbMy8aUYukRrL7ZOEnmVKX0u
3ZrwRwrvpZ2xDTlfko1t2/BxmkCrIb3+QpRzyDOcm2Y+BN/FaRRunNebG2xAdNNo
476yj43lHjUCiyqmpKa4HxVUYVGnUUx/2EasDIFjubzSn1YNir0I4hh2QIV6K+Aj
j3z/In68dAYlsdkK/RDAazV6RzSWQ0XD9wTS8OAjVPaCJQUWKwgMc4NwaECZSWs/
hkH1TfhEjIFjQph63S8rp+lYi1zNY2RiS9/3YIpY5A0jMVJtNVKHXv59K0jzVf2c
mb/TF0ht3WywSwKCSZ3jwBPescUJMNkNnLLipX5AOlMNdRX4Uc/28tWJOdpEKppM
aVgNDF0nrFvqruqpT7wXg5KCgGRHYsHUtoEvtySqRJIJzRENuK273Fksmrssb6eH
+D0iwSGU6hk324DP0ZR7jfGboBcEXrXoP89KMZlzIYGOtp3N/ScH644OmjnbnP8d
d9YtIPlldON+WQkhIygDy8KPMHFIKWksp0gLuLIj1pxxbAiaOs+75IHlFHi0bBzf
lhX1W3Fa7wTot1qaHbyYpHpUQi+iJpypEBF4x+ljWWmuSjgNFXGMsQjnb4j0YEuN
Opace9R+NRT77NlJ+ICSuBb8E0q3K56gICseJbDgas5V0445t8iTjz157mi5VcPC
hEAp6sSjS6rGTYvvP7vxd5s28+tAiYzfivn99kBOgLAscglHRkknPs5u79aKy7Pn
tHD4ovfFlLD1rggx6Ui9rmkOOlgWQS8k294wdBsYgPy+zBuzKw8rkGLDtvsBnwDE
90whGVFM+Qa1WLC61mVmdYgWpeo+0W8AyfbHUvIOcIEzNH/xgXghCQ/2TlyOmsPM
CQIXZ7Y623TxA8zsQiEwgiYOt5WyBv7CcXZSmacVMiaHLYrxmciDk3xJOAL64r0R
Plsc3PEjmDNpjrfQ7ennABMzbMZhJoEJu6GvdSyfyKil4LC+VuVdTDBCz9YykNTv
3piQfVieUfplsXfVnqOfOGddDIH1RM1plDHoPqcQosyosB5Rb70DOyyml2QP5VFh
wgpl1Z0nxNvdbYUORgSQkRVJ6NjXKPThlCCbbh+K2doqtrD/dSNzk8kClxHBm6ku
jiAz/2NypTNJ/m4aQv4sAaIntUI3Kl1/SmFq64Ddp4Ci0w7VJe1iwlJOa6tNXSvO
Lvq2KEcwJYZ1qg5dkZlc69Zybes5Y+f5KVib6n5O+1jaQ465sGTkSbRDQ4g2T7Mr
tiZF8awzcJEStkUjGZPFcXolqlGZCAEhIUN/susuq7v/beZRRHJ5n6YHf87zfmrS
eiM0IEJ/9zgFwIkfa/FZyUO9GFgXRGu4/opegh+7UEKof5RM3vJ/XCtBr1XyC9kJ
xVCsPmM1iXMPry4MoaXzeLrlH7y6EhWkTyKjT7QD9aCIUi8Wb3nIoHsu+rUCe5Oc
l93EnbF7cyBp3RCiGmb2dmGGgPQ3afv4JWkbOYemGJJogHo0bH0PBbAMQjgcE+4W
XTK/usocxevrBwWBI8RdBszMR49xTjjDPzCGLlQAhzXL6sb2Q0DQf0xcZTYr4D89
/0R65d+I0DhFaA8USbRbzuzmJYyv84K36aHgIys/mGj+m9Me4HTraWNykgbIpTOv
aXkVOVtHcVKDAa9dBoZ+mHa3oGQaAKvybEVvWYcX2GLx7a5La0ndfs4ihjLFfVSp
cpcRiYdx4R7ZV9SKUa5DQnp7zHsqjPbQHKacQfMOcf31vsYgDwtmE0+x7NtDUuhg
mo7zsqsmUhFXmMl4NL1TQwKcGKsy+b7QKZWnJ69Nwn7sdlOLSUuwnvgSfQIyp6Jh
VNHTNxekCpukrH8rdm6a70ah4foFS9j4VPjx1BzhExLTk0Biz3k3rKk9+NKR7IsE
BpkFiCwrEsYStlYdPSqgBDHq0KZpTwE7HDyqJDcQrdXzqZS6jwdoPVGqXJLeKQ4n
ITGxqaHyRXTpZ3TJlIPheqm27RPS0FOX7RTP0OFFW1dadj0Q3FnqS7B7NBSQUCA4
mdSyipax+ov/3KFrmSkvRJpV6cu3e8lVPHht9E8OfSNYxsbi1rKxMh0LndhO26ow
igREgVNaGEZWIXiAaN9sTR86leIvMIp/EznEVgXCw3if8ZcSr1qQ39LIuS6jF0A7
JrOnX6V+nQ5VvBFOuUTt2rSwNaLAmcaKUBRkv8sKZgNqUdqKgRAyQh1RWVpl/y8t
/5OYO3qYKqLyBNcxB6F3jmsr6Vm/uA7s8YAqxu1g+CUQSG7RTYmUvVFE58D58n0V
LgadhBcN+VltxaOVREWAllmsv3PX12Cexys+2jS8V2ylYZehIAaud/KfY6rMdme3
v5qK6FWRgfekJUA7d+uxMUkbzsnRCv/gbdpygsiuqKAFekme3Mz8BBg0Cyb+ZsD/
D40S7XMYX9UcNng5y6hWyobVpfDe4I7K93UsxJu+J/WK2h5aK8qoujqv2MwqLJn4
A7uMagpWAq90c1D2ipD3MQuXck+ZgTEwwUdsZLMLT9sAAmzPYPu7KAGQKlXmp4i6
B/JYgUun9Gk+QdoTSztPVr/v/a7GizgVOuYsS/JiQHEmq2WRHPR4EUiSiJunBP9N
A8GvFgORsuvkV8tw66Nhe40EevRE0ZfjeKm7X+4dAUlK/KZYlQ3Hvol9pedV1CCI
ijLVz+GBrpmbxkkEjYZRoKHFb2XT9pnTL+kCogmR/vqXVY6WMa8TXWQDIA+BWj6o
7JncCie4hFOCyo9SjpchyrJDFBKDaf5HTYsqOATmy7S/pxx1MM86RSkn6x/VQLFt
67uvUz5HnyN8zgAJMnZbJz2qbYJdDw7KBWAhO+GsCe8v4UwWE00WRzsQMrM8UkL/
GM8lQhoj7dJRgvmpgt7fY9cXt/Oiu3iQ5pArJ9ND7CyooL2fkFY7ax5rKPx2pJ6b
NFTom1gq4NpBBD3LN1aFnubcwAVJWkt5n7PdYuxU16DUOvUkYb+S4INoXH/M6gfd
8RMUEtwobPKpke+YIibzYl/xCXAK2tLGndHIUaox4IvGMHT1N94KtQy+hPN2DmZB
O9yLAfXpc4BThjPRmEFVvk3fEDo4cjyoQp4bHQhdp3/Lhxra1bGmsZGV6Lcn/HYo
FiCIE7+Sm8Lo5s6tbKBmk4Rdy4K1hh4P8wJ+4/8EQ7X0XG1EhfPvN5HsTrID3wqA
z+yDSinkhyzQ7jbCTmiUIwHasDi48liog0yKG1gJIsixsiraBdqfv+Grdvg57Sot
EUR69zd+Tq5jq1nnjXAuPWdXoLhS/d3I9qDTrI2dVaRnqQSFiWcXst5ghihmik7k
OmV7JdxuPWU9eVuh6NE+SiSBEcE02EwUUoRw3zP0h18kjeF8AqOq0NPqxEzVBsQ+
5xm6uHZUJOO4W0ZnZTOEMV9rmYGOyhT2StWk0nT4U8nu0+JCkckQqItoS/VjI+wQ
m0oTRWg8Hvtm6C4Zc7Vj4BZ38OEO5OpZ8QSQoXRSXeGgNpphJ9Qa7130ztahem4B
r9/EV8xncgJIxDysFe1ftYyd3WS9Oo9nPD/ZE7EFn4c6aOC1vSpTfbkx3NyhVX7X
bL56MolL8Vpmto7rzFqbtU9kiZLIc5h9KaUZCKc02JG7nk7y8HvGteJCQVcHvjGa
i81Ew9T7aJEFdJXHRTiZr3cSQefZbD+gVcSEeSi0kOyg5IDvHqlo/gOnKqY1q1JZ
7qiVXiMaGpV7noAM+H7mRsEdOBBj5rHozEAl53hB8aDTL3OZEb9NDLrKBzm5RNO3
MlPAEwNuLGkg8SHXOoKRaP3+a/bKJl94v8HrCstuRwUyDxH+aVoApOZMot0OlOMb
Os+MhXJvmGpub0/r6DIb+AXpfLRSSCXkDySPyFbSyMDNgunBN7bvpGuP+8DeyCeS
eNQXZ2Av/4WrLRyXrLU7nxBy7LI0B0xOOTcKKOmkQNJDS8/5ph1MRj0KZlTvplzV
98T39yFlQMM/ZoE8ON+779p2QIhBVoQBEjI4fnf2VvJ5f0wP9SDaMabwARfufU2d
fu7sa9ImM1Af17+q498tP5yqIAUFmjFvFPuQhJx4p7zsblwGHwyhtHnVPz3MK2jV
5Of2m9NjiZn+kxJOtWdsJcL4E0OsgPaKeBc0GtSHRhPxtixZHhRstRAgEARRzWRR
MLDMHL2ubF0+1ysgSib/Dw4vugsNOXF04yGmbr8OVEHgr3JFR7pBotyrFYIWVNc4
6Y+7Q9ytoWk6M8BvShq72a6hQpsuet1EXUDi177e31xscVC7pYGImgAbD7asJL2n
WZEDjr77AcqXx0qtAXR4fy8NJpXl+fvzuX1Z2SqOU8A/hdPw06p0Ia4h4jYvbn0M
NXySSd+c33RUbghhdw0qWBZ2rKaj3zm3eWeSDP22kYKxFAj9+22YbBQDZksiqC0s
DdjONxkXDtoLCWGqsAz/B7XKcE5VBdm+WPMfiWbSz1j2UFol28j0hDXGX+Qw/1+6
BCUbdzZDBiRfHxnLDEaKKNopKb4Zp7iEUXCi9C9keZijWg9u4tspQxAUNzTaSsyy
enL742bAGuEkSrTYh5vyTVkfHM31CXY6V6NSHO7Y1Da1pxVZU3kJDNxtFfaeO8jL
L1ptHppF4iJGGxwluGXruDfUfclnG+jFwgfHE+gakvlPF9/sESL6SAb0cNegu19J
G9dJnYOrn1RiXZXZ5hjUFDIMzv74+bGWYXo/uHwGPKEWLHEBrQadc7CvE7evDqXZ
tgkGwnkl4AjzqTOqPm6zzAT6Iv5SI9ZOTbeD5fP9BnML6JjCG4hXUYil4cIKPRf9
ON1DgaA5+s89Kv/ck7BVdBsDyK8EYy+UQm/kk6q9QqXvlsR+zPqjh83w1gnYMihe
x9Tqbew5voygpSn3c1Qd0rGtbC45/6z0Dz92PxPigp1WtxTGq7BWLctYsqF5n3vv
jDWBGTiJZUKJP4k4VlLUPj9wSOZ8yFf5/25/QQQQnY3OOojItII6P4L+uip8D3d+
etH07flvTR9RQH/GHcFKIhLzEUNXBQq7bi+XACPh+aPS368b9yTxgQS7QduQKQ9Z
tOc4fYVc04Cc+6pOPYBLpngiPYCSDgz/CMtE15s2bZof5efLSN3T4GDZq21fiPH9
QeZayPUbiTRBa23SWCLTYW3ur/BGKH8k66g0oGB9P5rZjn0LwzaLeGWNZypVvWai
n0kNe1hmvjAQr72BBU3tbiL6r+2ASIfAEb/lW5GEui79fjFNcWHO93QexB37F0Xu
BvtGG6JtsGzQL0rzXL0ybw==
`pragma protect end_protected
