// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:20 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gcehmMJWFcCLmfuQl5tQ6ZboPqAjxoYMxyvgct2D1FxZCgPijvwC/dOSyRquqKSA
VAf+jpb3dI11hWd5Jb49lm9QuA2bPk7zMcN42fohKp1vsOtLW0gDg7QDLBfAFNjy
XqZFUdClV4wYXMiGKIu6FPFtDQYuY9b364QVaqA8TMI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
mH17iW44F+eXZU6NE0vtDSFKUbEyujLrOftQP4ojbKZICIi6e6BqivZWNvLlvuZf
sgE7M4h7QGI2C1gkRncr+qlhVl44TAASYrkmw6p6+YGPfC9zVW+jCRVyZ6uYYmmM
jDuzXm/8TjmRfyZh+vbkjHZ0DJNyMg9xbt21vorQrF3SsRDy2d89mDOF09t4rIqC
P/k+67VFOjPAqu5oi7FmA1M0Eo+lbdkTOjugjhbhU1lWpaBrvrh04NAc3Kg/WkUm
aJjprYqZFTVjSSw9SA/nWsF9DgtxWBB5H3bDoPBKgTY41DYNag7nekM7uTNLPDlk
F+EOMt9mCyQLLvfcaDRl2WNr7LvpYxKD6ZW7Lk3rG9re0cG1AiK3zRjgPOlA8/C1
8UHEjlOOTa6njyuhiNuozs1YjqoDdyrIN/B4DqAZhrYzgIlvt8LHWDuhcdEUqUEV
yD1V33MD5dDLKzgt2aKUKQxW354adl/aySDeMOFqUPR7k3n0dvm0wNxqRX1VrT0O
axr93CC+MK51ActuzI00GBQuh8EKoJe/H2DcKOzKRU2M5OMbe3qq7F97uZW5ZyQ0
nHoKUbrF8ZAzzmdy9KItRYMV38raQpsxWKhrKL9dF/eHQUsKsP0eNSJKKn35VUob
vNXh44gz7gFAXq2ovPAsOkD1mIuQBShQvpKz9QbFBSw5LCKKQCDmgFOjeFfJ3/2P
EYZR0NfzuR9LG0qVEpflg3xEh8QzjaLVV7RbVa15LO6aL1DlgjTb2PfiVsoCzvZu
dAUHdhHBhtqagwK3R0NHQ70c9jj3M7fx7Wz5uUOg3Imgh3H2QaPcGZ/H9SgQE/pP
AfpwejrUyrZzghw+on1xWLmb072uxpd3lAxTYJLGQB1bVgSYpblBHIYgvA1qVhgC
r8ZtJrfmmumyDDf6Hlhu52SUXbhsSNUn6k8Ynk0v6oorPNUQcITnVQtTNo5AF6ie
f0LAIUA+KxjCeNV1TS94uS8+Y4frx+6bwTWJ/rG+xcte+zVd6ZXtttf5CcvOENcE
+Xj/t8XfRrajr8VlbClcoHY+sqkxzYg1EKnmGtNl+t7wvACBPWSonZa0B8f9cvVN
pNqucl5unNis38rcH2niYdrfCgN9zcWWyJ8t4KZTcn/+hZnbxAWqVi2GooxJoCsC
RFMMKmCt5M+twOVA6yOXIFaNJ+TYrryyWp878eZdX7I8R6J+D+PyOsRDqlWE8wpc
8MCY1uVl7gH5lqMdBE5lD6TgrJt+jEup99VjGUs2HaD/r5s/9lLiuIWx7/5ormXO
NB11+Es+YziqZXpkeyVv618ZnNw6HmFGD/QaLWwME2bv3QtiuUyIxu1i1Ffm0c7e
159YgL0b47NKD3HuAnz8C1n1be9vXb1TITA60rtyEaHEMf8uwCQG7lGChx6MFrFF
8y6+IrGD3n1of/UzbB7JvxogJgaWPOfjz6iFx41ns2rQkF0CU2KBFUW7u0zLZ782
CEn4epyNcMobODfWIAQbU1FcGTOm32PaKBHttPBlwbSBXman8gYgSg1Nrc7DmHzi
71OJak+PpgJjZScDfTaOuOelcwmdstfXAanX1j5Zlvz4g1wmgC4ZgW4TQXrsH28a
8ZES+KEltPtOJ5ct5m4P4W19yW+sn6K6GeBzNpQAu6vE7yrmlW/l2rFgDf1VOuMz
aoKf1WFSQIGKl1ThNm73uwKfR0OrKTqq4iUz1j1hjkb9vRMIPUs3AMGGzJZxoz9+
hc4vZioO2wh2PRsMnFKxknjo6jMxibMeg4tFUn96jNhUl36fNZ7wWfLi7bTN0rRy
+Ki+jNKpct5A1x7tur7tNhz/H1QFeS6gzwd5zfsqzl8giMPBHPg1CsoeN80UXvwK
Fm8j7TfOSLhYZTcL5du8Ukn5wep8BVYROohZLH3TjiI5zxzNZUWLkPJ6NZY5Cu1v
UVxMvi2xcu8bqqQzzmXk8qsTU0LX0JmF7du4frguN/a4T3dnvrXsluK2ZnZFEZgX
wvWL5WlpGcmIucHMChb9uYZBYv1AdRd9gymE3uXVp2xObWdgWiJVEX1xSCu1mZvt
3AzuZ15I5RtGSJ9pIKVCwES6vJ8ew9LBi31+9f/J54HwcWzN3BLlWbp7CVexu6Xy
Ui7exTFwgFaPnXt1hudKEzuWYuhdPaAB6DUlvUumy65ijVvmGwasFrkbM29Xrbos
knmd+6qv/1BKbhk/vpekgtd/wh2bQcPNx8MTkItD37G8t4OpzI9Xl7yKafnGE7GE
Ghw2vI2iY40spd1Kxdmh5+qbjwFR07O8CrmR7KYduwXBLPEP0/QIIHlbmrJCxHuH
40zNGedlECkQZCkNEqHExpqHJ/6LmDRKxEGQSzeFqGr2M6V9rOSc/Kbaae136PJB
+TaCSQhffPxMT3mzfhGjPv6E+2wyrHXjaOlyHFoSNLfCv4xUS2hkgCj9BiSL0Xv6
oWsHcOIXA0yPEy8vbawKjIBHotZpcGqjqs3EWKPAJoWovDl8u0MxaO9GiUEasO0M
fGtN46WqcwdaKiWTbwRZv8oZuNggIFdo0XHDH+ahYOjpGxOfxLSIn5C4YWa0llkm
7rLfVf4lhXMt/glv714eQDOPxYndooUA0Yk4XA3+Jz/i4FBKZM1axF1pT/IQpRG9
TUVpqavTA6YKeNhTT1UUsWCuR6ZJm+pRKPRax3gTVKJq+7QkgnMFFMhIJg1z9o2L
Lh1ATkHp4AmE71uAg7P+KuDw2s910/WpMou5tHfTbbNhKVh4LixL6in7RLivk3mU
keDrk3naXpP0iSunfLgUtsm8SQKQ9HaLJ8Z6Frv48ig+iaa1xEbszkSPeYeWbgCL
cum0jVOOENfkJ9rOF67rPhyZ5XinH/GEj41qB9cAfHTM2MpIjST+aIz88EyRM63N
W21+P76yAdieNcTXYGfaU54ErHASa9jg4sYZcblHpVCleZq51Dc6yHS7eh5YQ6dH
oSs76EH4Fe6HamngFresaSCrJunLWtx5h1KLpJOuY08d061YdJYMV5WrBT7XGHNK
cm3k9Zykj3josbBiOqwnOi8jTh8zXRy4ASpYW9lp1j7at/WJGfvRTDonfih6cfEz
mD6gBFxigvWNbXmKI+nI33wk8fCUQSP8cBq/50NwrKtuB7JaulULWuBW+M1ylCfb
8mLTq3ULHQy9Iqgfk56NeVt288D3EWP6ZtJdPgFyCZU0UOqKYGc2/2WIFo3kwat3
HXPxEbkVyUnB5bPA5z2wgh94h7Ag7BZVApaZNXRDAnrAhbSy3Jz3+0t4FYDWCfnk
0BeDI/XY6Vc5BH30NxwLBcgy/ZPYVTt2Z1IF+W3KNc0vhKZ684hlsDOASDvAEVKn
hoQvf0oubwNDUuK4Ooxwzl6C1bnETWfAHEVCiNa98cXtup6FnBf5CDXbhtkrXlSr
rH/ixF/pfqE7plLF0NuUrRJ2/+zU2Su/wsWaXQpYtgyeoMRxni/A/GQSwH2xOjIA
WK3A/fJwbTligBHpKhFc2yqQoQ9IvNcLrNcYkpWkaw++DDykqirnfZ0rVuDPzofx
HCO2bky5wQEoc+yOc4MYk7k2Nl/xODlGaQJL8MVUGU67uelCVYncH/wUckqdQ7vc
lPx13NC1CY6VfnqXcinxxSMxY14sePOk8IYWHi/V5lIVK3mgWTS+fNoPtQxUw3CA
qchF/xiuMoa57Z/AGtzHfxyWy32r2B0KTuARYf8PMBjdxKjVe9pa63ceCsrDyd+N
nIpPTFYaDaeUMNbc1C4pn7wGWXl6jYh8YWV1pjVtq547qPrXy6pNQbd5+Fe5Jcyh
8J+4UKgnPUAaYnBGIYLRuaDPx3RTLmKhavjyWMl1OdwX/RlYdgQF086Twgr2RaUv
QNAaNwYlW3sIObucPSsfy/UiBqoSjte9nQ7KlUyPHYGQWehkBmTjN9oNAYMTyXDL
ySNIpDiQE1RtUbpq8kiJvF5ARQW15HCEvhweePEh3QA+T5anFAN/4HZDP+kxd98f
TXY1CX7wZJiGjIc4J32hI74wFcYO6sxyiPMfAn0Kjw79qwpPk6PPAnHSvaTlzXFh
Gr/7fYLXPlbYJYQPpLMajjuBh3imXKvjEWln0SBQ7CEE6SXmkTqeP3Z8t1C8EywV
biALMxjzhfcdi8exo6DLUmscF4yLuipDPXh5iFw+jV+QPvlLTPWgo6x9tsr70TWq
XVR+NRw+zufbER+a8w3xjMe9slsqQR3WJIyJ4yl7WLOl4FgUR+jh6E63fn6fLzz7
IGw/+fk1qy8tZabMuz+T4wWXmw5oyN/q/d5bF+jFz2RooLIjSAkmVdT4cENtlDbS
zkxBC17eweBtgsjqYPObuD7yMq5j/kOeRcC6E+IsrgRiaEdj/ccLC25n4l6yNxhe
yjxj4pRDChtY2fNKd8/vvTYteJDo+r5nbTHldYolSGXFXvz37t7OQ1v6ezPPoKzA
Phv8REGUrdHeG0RgfF9OB1zkrNtQX8Pv+OfEqKgYWbl7oAkeUR/hqyLuthfv+YnR
z/AzVx32QYtPFEBjfHlKGn3DUjFZidB5doagsbWm1uNoZpSmYOcawPl0HQPKE5d+
KUJvTte0qmRwm/jRE+xuySSBwOBHT4pT1nhKbZxbs+jL1u6BABBPLMliAw1aL3vQ
70DUCj9Xb2hAQoIgseI6hPZYUdTwH+9DviSCGla0oAOoWMRGzh8iFOkXQvU3XG5r
m1f16Vw3vhJ0fW3nHkIHPlrEGZMz/yAEklM6JgbazSNDTvpurMnqTOUfcPyYT9pt
FhgcvVaugt0br0z+l9YA5tijQdXbHxj+FILMGYZdfr7f1MfYAdPwnbsPTL6BJMI2
YM3EYC2Cu7T49A4sUGxtDm4mtuY+bCP/lfJVEU09zZ1zUe9FYNsKgy3vt1sA8c+L
6iqx8R4zTYxA8RYf/tZPyUfaH/+Vzjz/i6NQGpgZB0ytHG5NlpSQLsXGYjtmV/O2
Gkm5WlX1Mj6cR5iYZG2/Z4g96EdlFN6VlGpgppierZ65h95gXe7zwVkO4wyyReqO
HpoA7YYAaoOL7RxPs0eVAYvbZSh3cJ/1WdKgs/Fwg2lAHnsvfrhfbFUwlRTw5Uhp
QMYoY7ODY/ySB+q0j+b+q9OkswLyOAgM+eF0+W27SDSA3BVHvRMlDTI4xFxRfsOG
frQ+pchU8OEtb/dP2iZ1zsZ4RwWvOGSyaHQQhrk6rJJwZixaYWfQsnyD693MwAC5
AR3IU50frrraYCOdOg0pknhlDjr0iSINvpfABd05ZIHDBMECshYt2+2bC5wGoXiX
YmRRvkeRex0RnRggAxGD109lgCrF0N0001DLxmLc7wNhvnWT9263/sZ9aaegRCAt
o0Orbkqvmm1aVhq9zy4Q0lXyBNH4HuSU0Q30r6Dpy+m2napyesyA4u1/t0SLispd
5MLLwRogNGNs/kTnsBZxOuUzOe5CY8mBmF6LH4a6VjN18C5WbCvF/o2yCgHrE8wz
lOB7Vffa46r+53pJr4uDYuM8cmTJTcmvtXSQZjnWDR/XjU317RGXwkjn3DFwnWLa
YDyOzoYhQdnVO2QeAxT4LcVWzt6qlVy5nCogzveUQbF6RVq6K+mqBZZkTNeCFSC9
qAU+7lVefFqdUk2vVOiPmPG2g1sfyto7fbhZgeRUhLrNN18yUxXW4bXTChpBn8c0
T1hcop3MofHqIHa3VuB5g9jIwFwX0hCtbLTgHY+OCc51UMIfSjwMIgBqQQhvjIDL
gQkQHJ1XiFPGIROHdlA9bCr8GEVX/J+dhM2eE0lYS6ck75A9iYuGYR/ksWYWzfLs
34YnZ9cUYT9uxjieXCaqARXQohflJFH60O3hkeNN7cqOftEcwVu4XCW+1mM3o/Mz
wexRxZCtiMQrH/ojVaL1KRrREeOSg5F7pMR205r8iPp27kMd5/J2F8y+HlUilnR8
wLdJDUolxyVylIV0BUVbUbAkHmBDbsnJ24bKAFTEEQhrLt5HqEf4xIbvqgQNIfs1
dptdS9SYK3JoziiGUKGEz5IOANTmmgbCqXsLoXG1SZLy5L8p6VIubGkxJyeZCbXh
nJkafyi9XPMOhzNZIHsHDCYtZxACu9HG7etoR5sLvSfLr0f1jxRE3UEw8BZm2dNF
9B7wAptVhK1zizPFwAF6P0zXs6mEAEFXpWtQV5QQo+P9fcRdGqY/xvteM0hOg1qK
DKDkHefetbz/+JoGfsgCVeqGNLW4PUv6Mius2dVv6FTwtMSjbon8QuqLbymIgQ/+
8ma63JUmFWQL7Sl1WpcSFYS4R/YdbkIoi0qMNaTaEQuPv0b8HF52g9u/+L5xdM7b
IccSzE42l5dKxyR9BVAm0kY9qYxBjhyU9pcvzpcpzi4iQimSLZcRoSrLXgC1KETK
s/ULcMyjDseQfiH6i8DNXwH+OAw+Y12wNYN92jbkyV4g8i8DBSpiMdppM2DejFU0
/s0H2baO7AQMcDQ9eTvfV4wH4Fyn5xHkE3qmQHqlBnlfdBD8XfV9rJ/6MAwAUUyI
0TvGxqZgrQNp99Mx0GpHAeo+1JiobGUK1dXSACvVCxjiG08c9v6e2sibUyWf1dKe
OPr12a6kuiGQFXv3x9TmsHVhi1GaKjMEU6d+Dk8GAJDbTRi2fxlyTQjHZcavIo7w
ROKwQrOPMfFATvaohFXAtR9NKOTRQJTPapjPUhEAgXSrGql2K7sg2goH+9XBiMRY
TM/SCn7IIMsIjZe+MavsYpYVWllsa6rzQBMFn14aDoEjWKZZP0RoU6kDp1E0SqKd
N+c0wv1vpIoQTc+s3bLtiJFLEHknT44obOfafHcybiA5ReqQGgkbRWsPrCcmmosv
3hK9YctbBk4E79hd8qa0Yw7r0446V4xI0VBPidx3m4LHCZlolQn7yFinuVP7QNWe
hCrDWon4bShByw3FBBNLzB3ViUwxI/ayv8yiX2aW9kGXglwC/d32nT8aohoc4s+6
uXYRV/ZtNMWqRHzUj+M1A1T7kZnFFBny+C1GBSiyfPDi8YByIRBpvKMhuQ/ITtp4
mxzaSoYbfge11CPSZ3z38GPWbK/f6ktZRpD0QjdUjHimCW2KJ4EIdU7g6emKANNc
tlxMVZWrn1f+gLe9gWIgpRZ3XJf9AsG3NHqphaYXtUvPTkOy/uVaAATjpqFlNEgG
XbZ78Ruj1eGJE1GiY84JI7dWRH2M+jdSb570OiYihUbJq1EaPRGfXFp/sa6n67/k
8XoANdbhZ5nZcv3gYZhohS4x5RnaU5t43Sc2OoGrM1W+e+UnMnd1s7gwLys0Sk7M
jMBOgn1vvQamSKVeFHGWNhvh5Z/QWNz6+WqNjxIlkTxdci6wJKmjfHGin8Sxtp3Y
vonYlc+nWgv1DH+R5Wq70PpEwVBgLbXdPhh34b66UyDvr8SuETnwtwEgbBpv4DKf
99b1vhjfbvJsZduclSRFCRlLiyx/8P6eY9EgzC6nJwcWAE9sRtpXpFLIbxdVWSzB
0e18KLcztiExysgWz9ZHUIzOlEFiD6B27tthASX/35ajLTx4xvFH/8kt1inBtrNg
twzEAauMnoFnah7DAG9OXbFn/axHxcNqTj6PxShOPnAO2muZcsEkexjODMdLBR6W
yzUMidjODpNnVBdyB6oRyW2zk2IhNBVrIkKGZWqY0h72C70Q/nafbGfVUjZfQNhe
ekSqq3pPoYiVZHrA4nitLw==
`pragma protect end_protected
