// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:15 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qriJQn7D0cwg2YbZvroLK35O+ld+DrAnHkgDi8w3NI6wNtgQMX8IYcABEdwc06C9
gaWlfABOYoaoKiILry6udc3LQEa3WKAqbMMq7VJyXEJRRGFf44dqcORMQ1Am+BPA
iPJUiUpSGf0ZyvyyLfGBAI7rel6lUsRi4aXkmZnximA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
BiN9K2oajLkFXMUgZ7jdVorgQlk30UMLVLx30ME9XEv3w2FDtQF8w/ykd3CeJWZU
rhTqCyBlGhD3ws/3EZsLxG7ZKEZM/F8SbvrWF1umNCglfp+at18hPp0A8eivjh1J
YZf0KCCUC3vyidVg70w09M0BURNLs1LQm4c9asG1MZS6Ax9l5+NQUEV48Qhcyex7
/iXF4vwSl9/U4aZLot70V1KkoBwgeKWNlrftCD1u3b23j18J+jHoVVlcHV8RHHTN
N9Aw2YCVhsoLOd7VJ3l1HSlXewCZ51Cu5RHoTj+AYxM23peWN/ZA62QTopkt0e54
cXtAZk2wYeEBTp3eXDZDuIJxfsI8qhckjOg9fdETdgn9b09WTfbkF0XjlfEYZ4aM
V7lBITJCst2I4XiGkgUUoaBW4PRk+JtiAwkujvCZeAsAuoR+wbEjr1Lf4OCZxZ7U
ng18kg/LX7xc5NoLwma+gO0/NsJOhDVvOZJNUUE2je0IysEEQsF69lsypbEljoa1
AGkgRm96/gsdG4Owk5xzN770k/S14RLNbDyflCbfh4cS0G/Ivab8NyBc3ofnf4vA
U7sF2ByXw1rmRBw711+QysJd2YtCrE53lzZ1sIGFbowIkc/hys9aoBtRNB9k0+jT
PKk1VSacWZ85d1ABB5bB8O4Oe7rDyrx2ZJOeUg7PxdnI6qp4bRtgXDJSdZpq27lK
0vh2enc2t6wEKIZ/Qa5cfZDNA2VdQx8QyJSE67YWNS9WMsTFWdu+BgsoAovC19uo
CABV9jDenq5IGJ2Q+u7TyifiTBsc57YfI4xHB3+BeDdXiyVpmvpvpSwkoSQ2OouO
TvnTrXy/CVVCtrsdZRAsI5keiwn4MsUNzF+4JHAwrhD2gddwoxGtzKI/zu8V/Gi9
I8OSsZGPtnmEK0i2KVcyNDLvS5wb5O+6WmMzoXMjUvRqgVzC9KtBw6n8MjtzIIJv
n3PIMkTX2CnzcsX/r8Aspd1f58NArWgk163FQFLbKmE8xAE8yz+YFHsoH8UXAPis
SxMwRUQCQUQztD3YAaFaE6Kpoj9mMqNLZbHTW4TnEx63POMDH3ttO+jNH4XOdlrU
ys/BdLHIeV/7SkJdR/k1FLA8fLasiWmg5r9wtFrk/0L4Wk6wO4sApxMbKgIaQWkt
siU3tDD0fMq4G8vwleVIlU7K1w/tJ4nYyYEroBVu8dDfAiIMrAtqTX/dGqRWHWOc
7EoM+I15THfA132Eb1O2NQW6w/eaNi8k764isHdvkGntSZKb7OKd7xvSuTtSmQ4C
gErqCnEmmyH9E+/5A8ah73dSkhVeYu6r7US4yOcTdGb2ZPsgJlyoN7BnliIQuLkN
QnSD9N48/H3ArFnSlxFa12U56C0tFzPGK0hNG1iKacYmwZpdj6gEqwZ48B+Vmyn5
dQ/rI3EAhIN1wPZsDgZj/I+UuOfv5LUj4Adv16g3uvgSARkTuTAxA1lPv1NAZNl7
BYBqxLj8vDYZhQh8TPwC4/w2OFM2bgAgbtSdK/aMOkPQAzCDJUoRxX6QyoVFk4AK
TKnrC9WbMMZS96LaSgjz+IV+m4ph1bnNvWtZelFUOm2j3HapKMUjdTpoRv7iJtTJ
Eq+P17TgDFPJq7/dFhVHs8L3z9nUv1skgIOdSoZhtB5sfAjoHNb4S6WEEOpNGarN
ASQf8oaC9ftU6cDuQmzscU9ZqoSU1f1xWbrXlzyYfmjKGkiPf7J37gDsg+NZEeWS
ppAgZhV4+0bzV8cGMrsMKwh1oujqXR0knRc1VKSfCwdUS2QFO1QSH0OSao+kOXW0
mqCkIcnByypjsmzGfecnxt2AX6aSmrMMWUEzz0CbbMOoODdR5MTnvYFrdCXy0U/P
fUlLfEeaCSi9MQn7n/IVwfyei7jzY46QP+86LaOtV18AFIPz8Ixiz/y0czVFhcDR
N0F6fRFyAesSWu1LbRsOFXltDC1p1nNR509ABmT2N0MpQ9j85vyNAWNXEaD84sHf
m3kmDT3rAxQka65hUTKkeMfcRBas6raf1iYHbiA59m9SML3sNSJf5MgrsIXIOO6i
jw+A+nNnrHmLzkXsa0Qee/WkWCVOGxGEFOMmRksyHOPtQF5bS/oVKNxXGiTSdoyc
iG+4ojLCwus9tZNCXOT+g7uxxW5QY/fcEk70KYKsoKCdDqGuc+XBLOH5TKxXKzoi
PrBLaDuQLke90xRfpdcTE/iIzGfm5iiCZ/T6RuBJqXS3zIzlOHNZZ9p5xCT9nr+n
QvmkNmzImGWxdrf16I49f2raQAAIaqhZap4bdw0Y7GuDN8ZnTj3hczDVRFCq7EkU
UP0cmWcuJ0AtgM6GYsECwRQvxEm8BSRBmYcIpz/kyBt4eEtEpKDaLRYoUYqTgc5m
kDYd5UsibzevOPZBUG8w/SpfhP68WekyOi6G0lwclKTUyb5o7QvbcAAgqNoKnKuZ
SySqm1c9v7PTpBey6hViSe5UfYWWkv4GPsSoEt3DPyLIUoEeMsaiGaeEkCgKDhBz
CV5IFfEYjhfWH7DBpbhSJTIJOLlkaIeBXMpjgD4orpxhhnQ4x/6AreZokfNI1yy+
063j7m6rq6o3nZ7u9Miz8sHbCwfieffOhytyDYqkNzub0eoXMhTMrVTSB/pYVQNr
WIqrvzMKpyFdl0IUwwWc+eHpjCkcp2MnptOTpWGMf/dkaK1nbVe808ePBncr4TcJ
PVWNgA46p0b+2JrVF7hVEpsKDRWQY+o7dVx7MvfBI7KntOELBTq/d+dopPff/3oI
Jkxn7+qRl4cPjSMY1i3oWB6k52n0erbBd62HKm2Y+EonyvnmjOaFdxtCajXU8R/w
hH/8nnJH69HKFcXiiJ1FBDrjNFCmkIHFB+ROS/3CKhtz0e6f0QlZYIKFQpGt2Ogr
J3CGLKaTb3EM2Z9ntavF9HXAePOoqDZbD4myZeJaqINDXDudBhiT1/SZT3D3bQ/+
OvYyVo9gZ1jnL1c7/cP/STfeZ8JP+6CPOqE1gqFeKq4fz3bd5K+Tu0vhwDHj6j8G
pt1HAu3Q9yn01UzXDpxRCBWOWIA8fFJnM5C9W8ngJwSkWrmyxRmkoIDoxOCL686l
kDLzQixxAHrzQNl1cij9WjfmLup1gPis+d8iQNEjUDVdChEydak7PHsfc1TA9pvu
dmAEGKBNArjTEA8VddEOYCQXYRkVrcAzkY2V90IqE+VFGPbHAbLeg3Bew4fiM0Q5
3sqj7xxWrRbsUbW+SaiXUEkDf+fLUL9lv5fjphaO35pXJR1clwTp/0L4cmTDzCJK
iCaGRodU1q5LTJBwO6M0HAVBn0ZLIY7XePvEGVJ+hWOOzTlWGyixij0qbIIC9w4t
o0YzOB1Pg5LJ9Ku0oa1T7SRHUBkK2aavyIVzR469HSVKgsDR6wLl6a7mmvj74uk1
BO5/yhAylb2xGYhSnR1evLhT2UKcYNv9vH2rheKPLShXJgwd9M7mo5+zPf8WbUh1
Bh1IX62/JKyCYRgWeBhzB8ro+Adq7Ue6c0Yygh6D+P6Wlz/EHuurAchSXz+qGB7j
ZR7cUppcLjqqjoH+RyZIH6NftcD46F9OfG6jwPTbIf7ANPf0stfrss+MuFHS3tWt
ASQeUfEiVjkj0jCaOrBJI/y7NV0Ej9jlwrl07vDp3D6/SZayGBSvzM632Qtq8oWl
b98U1ldZ1ttko86paaRZ4w0aexRhfHs4NXuRWMFNLQOQR/8erTa5EGn0TajebVVF
j7opGQ5zt2pVSoaIyUdyuzcJS0Z+cTXm3UdhUMKHtq+YyXmletjnLkFyxwTlFkUW
ln9ztIs15WBZB+WlwiZAcT5rvux2JrHPSktduo5jYrarNawOm+P4DS4a7ONy95XX
PmvoqTRIkpjaBcNMYDQTQnd1/mbIQQghlzTGBTsVeOKIQjfXPBJO8UrQCUyLvdPQ
t/RB5Xq8yFZSuC7PfXCOMutroKNDlifFsn9ARER/fJrotbVzAfhWVQce77rhsh1a
uYvE9t79WBlmcFOApBN77xJdtMVF5aEcn33BF00ZlL7aa2VQlpsnr76pWTITsNkw
iNbloiXeYKG5xJ4SnSmFdhGMtKHxFgavFkKJNNnCpWzozbQKy2Fz2YH+YqR+4fzV
3zCFIzsfYy/SeweT5NcTwyA277gYx0GtjkCgr8/+4idSbmZaxz0RY02CNY+Gtz+C
FpQTt5SxVurio5PKR1xIXliWZdKWGeebc3KVD9X9HfBnCgnb2wCVMo4FyavQGSV/
RHKUY6TOeQT4sIB2LhwK3aERlopmP4IqatYjw/jAL2EOk+96c4hGa9+Zag/LXiId
bEGRiXscYHLrNkpZMWeR3NaKTYtnA2GbjrAwuws7qHbOyPJ2eWAHozC7srqjo/ZH
LT6S/ZYZK54e76vMSBY58XTLcqEjoq9LzJkID7rRUBFnpdt74Ql5dPI0xLBSmb4R
wHveOkJCHEfvBht1lAswsyxgoQ3nY+5d+AYY9P9tYt8V1OGQopVrAjokLwvLwNz1
hxA4LRw8TsFYC36Y1zHtTVQbwttitYMxwoblAUhxIBrgfU1EDlLFb7DUfTuioCbJ
T60SxMz87IX5TbzQWeDWcevdJwmbwWy/Bs728l9wXyZUxgKU/Hf4TGR6qPKkxAKc
5R/JmTf3r49bX2q1kvttUYL/IXyqawxkBNK6LcTcEIeg9emalUZiHg1gBeUtGhmw
ENEY5pqRslXyMzdXa7Cvb9U4AGHCG4VHfrg2ils8h+IAZi/g4xhgGoFUek7yu5Zd
p8OVlttDYFgdlAZqiB3VBOxdz5p3osGvjXobz4Ga65UA+6DUPLxd9g0RiIBxQ8Lz
yxnZSV9+42rjUoeLkaqSTGBZFq8/yFvSH3raFGcCZOyeyshAM4qEwZ7mIeo8cnKY
hF3Z9JPwphaqjgOwtZF1+X8SPZAFEVNFzvbaqHe5kQv8XbyHhoQGZ9zwkjiuNry4
1aRnfir6aLh7hfPOciWoCqcd1YO439RkVW8FExSiEB+ANFAg9wCqac4IrkCIVWTM
0BnWDy55DU2YUrINx0qHujwhmgvhJc444DFa1ZML2s6ziGeGnqfrHEddIJ2J9Zv5
cH5o/lCKUdwM2AJjBU756xLwweCZeh+c+gm4PeRUi0VyXAjn0SkRM1hHPnJIi5T+
zjFv5FHOFvopEFrhrYvP22bCg+FfOAPW1xB37YPJBHlWqMerkEJaSmAo7734byvV
YK+/pziKteUkorCwpbPc5eUgnvf0n8yZOPum3UXPvK8bIXVIIt/bTHPgxdbofi2q
2BdQTUzOg2JTmedwN88feHY5+5tBEdebE65yx+c0EL/8DietiJ5z4hm1J1Oqa83Z
gBSz7a0vjNtX6GPWXr4Db1C9DpPP29hDMw4xuibdGYybclcfHpyV7nEhZ3vu2Fe5
/WU/kDUXVlRAN5fAy5Wh8LbXWpb+Xr0bzlkTaqIZsS7SQ4XJQW6N+qGTIUYpR7n7
jUVQ36j9MU1S+61avc+qOeT9Fbx1uMRTyj8N0HfnVdbwx/+QuSdkfJbTWaE1Uj3j
Wh641EXu1HsYMNGblcm8Km6S+fLsvqz83abu3VHA64qgmqf72J2oraSaNhwpsNIV
ojaJOsZIu7pctsWkiYR5Ov6Ab0trURbdNUGpx8zmDrCYZ0RIZxn7f4C1U6KXgg4u
74MoWQ/+NFm+MPpDkYtCj7C0o0q1ZdozlEEnc1x3Esv33nbYfGmP9nvUYRuTfKSh
8NUWhpbqOoAp97VTm7HWVGzNxLjGmqAI4e1Fs+2EYexju4TcHDepucKYflDYVZwI
tUTWrRkqt0pSjFVcayU2meUndjV+0ApjEG6MiX5QZU1L7148W5QB7zP4nW4cLdlm
Eeznpj7weqpafA9RXq1yIpqdTqY80rUWHpZNJoY4yki/X3C01IgAeGaz19QI8kJ3
DIrHQfjGSc/MZjihI9tUHz6rq27TrrIJObn+H43Vwt9EoafPThA5hTa+Bad/qNAG
NTP4SwHesrQPbc9In1798FjHRLIHrPYoRZN2bs8G6U5Ln6YZYB0btqSdauRdHxhi
PkZLzOh/2d6F7ia/QmYYFQEac/AhsuT/xvbaxmSAJA47rfEqRwbaxgUwNna/RmSO
WyLL4Lus+fdqExYVVFtJiyORXtV08eYxi4Ic1519xI3DANPE/8IOGYyPLvAARbBH
svPdto3oY8FVqgvGW9crm7jc+BCoMVwedamYQAq09vjMuCFF1qPoIPshw0l3TeQ2
HC9W4e8IGPSA3/gHOGzGO4RBQtRTyCPoMaEGIchx1j+E6lgFzU1Uu3dm3rGYdH38
+zehe7BBhoNzMXKa44XmhzRbD5BqvhD7VwsDRTv3QUJ7PNYUvLsT5dYXjoemhs9F
33syWPrEV3aWZDoxudmjUoQixhnBplyLWG+6x994XcZVVDLHlg//2ZkLOxFVv+5n
64cAN08FfMQ1hi5fc+QHddAXkngF/hWJX60PWe0Mt2H4rH9APAiXxILV/oXGA1d6
8ZVSFiKZSvwZxzrFE3L1YJ70QPAz08JhtUJtdE09JPm8yGAP1pcOK7VnoHlOmUDX
YEfpNZer61gG44HOHjhjo8CmYwJ6jOdj9zJAxlx+iL9NO3YfMnDBxU6GVFdY3E7v
SzUCLhtKEFpdsvl7pRlG91eOXCHKibFLlVmzs4y5abFdadFVbpCE5SwaebHdkXwB
XIb6+O00Ny+VlrqOH+WeLnsjm5tJLk2mA90LIV+CXS5tWl4YijV7zsldJpTaXSpr
cwMS5gPQ5KPvI5SJ+IVRBqyPGm9agJHgMKvNJm9MEKfB+NgPPsvaAm8Vi0nXYPH5
g9ojgAwRf1lJuQkHHk5TnJXyj+7cgyWKNAPeQeNrFoj/9o/7hkfLD+gbMk7EE4Tc
TRDob89JFjD7sLAM+k1jLatP2DLufL20aDTjpihXBm9W0gwWzIAMaMqwj+wA9Rbp
1ZnclfHQ3xhr/VbV3yWf+Q8Pb7u9L/snYTGhvDbHG8xc2iQ2RCETWuLHEqOcLdsi
26f5LyjgD3NlG7Tgz3VPl10zE+kKj71qsGI97lOoxkyIqghGsmUnHFYsLGNbPjxf
Qm4hbSeWmFmpo4Pobnowf1TZkBcjSVq6ktIGwtzmQ2iY+hVQ/iwYn/cOYF3PFfiE
HLMgx3eOOrDchyl49Y9yDqLo9KeK9KHFqYJTWccFTBXHaJDXe1D/5YLPADxiLSbN
pjSPcTRplJs7azJCY6iKSfb2qJdbzqRRhHcOlLECcnNP43bZkXRHhBP9sQ5Ts/hu
7ih+QpWfzz7SVk99AHiodkDwXxk6+NXODdy9spVbL38iaZFxW8wQVTS5sjmvDoQy
ZJzIjdgF4EfuUFmQGmtf2rRhjSYx8ZzfrnIUHgtxx70KNN4a7h0Q1kfZBPoAmKU7
FGhrWjZtXF4acxa+At+edWDPHesyCSJ/Uv9nHHAlomuD1wdWj1y4xTrobKuBbLC0
h6gzWuEvEV1y1UDuQZ5amZntJX9gD19sLVltp5Zcoq+JUYbFDydSrHVGMSfbNM5g
XTiVxiGSNEtwiQLon1qXdlUXi7w+wgSRpMrsApiJKsble0W5RVo79eP9Zst8AhIV
GNNByBSwUTT0vleny8OkSpENKUT0qYHC75HfBpTKaYStl4YCorjWwDqxcrjl7Wzf
bVjvl83ksvh4P5TEV4IqpG4H9/gNja93Av/0BJa2adlhRfalw7AwzYnyTDwSnIMb
Eftq+957e748Fm29DkdvaoRFD5MjyBltyVOr+pk38inYxvbLzn0O/ScMRY8wIB4/
CqcoVT3MYhGKr2SfZh7IrT/HwlwXyGXaGUxCJMDazXWNRdyVDfhASGqe/gY7D97v
yopbA35VZ2RMKwMELWthl/1rn1uvjW7MDmjSwdZI2rF17meirpbVntVZjMPYZbBH
CkHBRZot4QNAxrd80JqK7//Z5jvhDAb9C3U5TwkcKG6lg5mrUabx6MqltkPsfr2O
swMK7rc/dazb5PqyZPx6bZSIC2mVY7MMiqr3faRR27nwN7q3yktMXxSrf+gfAVHl
yWoly/jYkLf5J7O/Z7UFSc9jbUU+9ZQ9scYeG+/u6WK9tlQJWWp55jcoU5FhM5ND
mL+g7L8yDgCZIhGaONcSgzgyvMC/ekA1ztODQm/SNAdcHdqHD0ZTjqK+kpjhq+Jd
Zb1UqYfUkGaSM465KtPUBFJzwuOSwdicmq6+jrDDQVeumv1aUPBCmqgFQxlV9R0i
e7fjqAgJ1+k7iL6H4Rd1hdbKlkJcDFW1DBjkOZKLdARVNcRLP6uOf2AIKuipXZJ2
rSWZKI9/RYD+byj8Xk3o+C48WGKU3ZzAs518LLkC+cZUrVKI04z4WAORYUJrMvpC
GrGkju9Gwn02QF8ZOBdrHU8g2w8SAmojZsFFLU7sCc7vAZamzAPatrqwpw5EX1B7
+1pQDG8/3fws1rHLcnJ5iIlVgBxbhNXVQE2LdsCHSwxreORjvJSnXreIcN9u0PY8
7zNajEAEeQuySrHt0JvV8kwmc29zOYVTi+ZGfAdYtz7N4xccw3MY2+9uUe7kwsQp
Msy4Zqqsp45T9o5SXyyiLeNzKMDShyH6Z7My1sCbLc24iKcgXSVPx7qkUixCzNSP
2Bxbi87S4Fenc4ZsiwCBDqGX8LJrtA3OnAjbirJZJYEA9QXvj0XSTuDkUUg8qHPg
RqqiAyddna0mD9AxkTMQDnkF+1V4z+yJMoX5TAZpj/LTrbKw5IKLNYuVXl8B8Dkl
wAK4T0KXf+2jHPniJx1H6+aCiD9lMQM4hLvKrUPIzIgXtKu5n4PNO7JP3+y2cHRn
fwWn6fwRNFFXxg8NloNDApqYPu1RBwskY2jd3YwQ060ctOyR5D75kiZ/G7ioPKL6
bijDi8RIpuKGSwdmSOs72tiZoRl7Mla9APAplfgX0AEnBCox6nVk1dU0PCCHkBRG
4oQLAhq1TVX3icNCPXIkBZZ8/snF1cp/ktyXMtnFswDl7S+ZH+Wexnun+Kg4vQBl
J9q6Qgl1tF9unDhNADaLsZlFNR5epVujPlOj3qlq5GJ70ucr16sS/eH6T4Lrivy/
nAPgVOuYeL+wHlPo5/FDvuqEGTdUJruaSQY9JqrcnRvf+hSnkb7aWbWoLI8OPskg
1T6IxlnxQF/6PBKnuv/RhlHZfX6IosxjE16djuhbq+nCDpPBVB3cgpfUiilYBNdP
JrbBSjgdaqFLHORWlB6OnJ4L91ilHRPEpmgUAHDbxMko7IeKnVmEQ+SR8xu1wWBh
scTafHHNYNorF385uBXID4oMYRrh+AqLKjExz6NTqYKX6L3fbH4RE/l3Y1yvGeLs
nQkXeYBJvFIth2ETuRsx/Wb38eV/7uOspfWw3a7Nyg1pw3yr2EDSXkKST3GRtFHd
4XzyQOQQ6diyxq6mB4TuhiA9OD/I/PjX5e9a0FXJxmv6M0Qqem2oNy325Ph4dgLr
aaG+9DIbVPgCAH433jJ7uMc+NifMM/g+toeyQW8gshidzj8ybsYzC7iwnsT20DYM
9oT1XdT/s5ueKQtDiHFCxs0OiGYAtsmj2Yf8sicwXu9En7A53av2EcmFnL4bUxy0
vxEjLVzZv8moGfLUv7HgSawn2LS3rHzcz9rsF3X5a/TBxe8v/52FeZ4UJbvk50Pa
8NZRpha0WODO4uk7j7Jnc1utF3OQg8P2hv9ZxCWPMCxxMXrhACHKO2KrrfDRNS4y
vkSjPWEnfOrxoyug6y6ub6q+5nYeWE46B4lTy2A0RgC08mva1Da+K7u45scQnU39
3QlS5sodD4orXmG1ZVzzxQg37ujaLOfysAF1M3mKMhslmNEtyy8i3wJuS3XOBeOa
Dh5h5UyUjFwv5jqoDxyr+upiS6krrMC1ACu+pUBjRBXBxuzaPvnAwL5I2leJ+aMk
ZV1D1td+aSCqcaEV+xXZmcHLs5PkkT190ESSQI8nyh3JOSa5ZhXqW9GNkXG7DgrO
1d01SZqgbu3tMlJeZE2E1RJ9L5VPwH0cRmQLGT3YsqLmFdOzgZOvh4s2n9Lww0r0
a/c2N38/Oc/YMK07vV6swuZAIbc2q0WKu2tki4ZtvpjBahPbzS+ADpDC3GLpfDwj
0oHGpGWt6g+E2eZiz/0GPpQ/EGbs7PvC2E9qDLUGihpKfZLMKmFXeu9SdWrbpTtS
78WRLbIqB8OVHg8vUmR39CJDioVcoWe8UdFv1AZ/9nvYB7gIGWJxnPfs5v8nWysn
u7uIz4JZcFKLOOcfvMJCzNoJBwSB8uQ2UC45Cv21jCaPP4pi+4sdSDvFMqphoFvC
Ar68UwP6G8YtqfJXbfkw1WnL8/mqWBr1eYgImBKmY3deBzn3S3KDlE1soSmWPeF0
R6EVWpL5ywLuA+2vv0sX4udzP0bLOIduSlmnJr5bO3hduqiCaBwIFujD4PL8XaBb
sIMJLR4ptWUM1wbC0ERjxmJB8ZK+mbuPBGkz/LAma/uUytryBm4psp/GSun4LRqx
ibNaWqTBF6pO2AnCyiBiwCxUnlbCXPBgbt6qJLP3PmdOpcjDx8L3m/Ci6J8HTS98
rltm5IamoQ5vTx4TRUSoe9IsAL79ou3MtAHen0L5kop9dnMQsJhOAVnVWc8wY4HE
c5yzN6VTPBxYjs9lQg6wpLF2hVt35+VDN+DMQ3nsm8FczVRWC54Z+M4kPmuTyFyH
LIgi5cNZ0EgyZezejISvAwQmGtkYY+k6ROaxxeycU4u530eKKNnp/66afng7edAZ
GfrR3R94bjcMvTgG4zOJeqLr1HXZdXTOEo/wVeFkYmG4cyPGiGbxki6GDGKFdG6+
5OULlOVrS/AOV8/ZFf5dSz/1zf0EhDakuHi98TGkQ09wYLai61vNlAkNq7C8SG/T
at0Yau1rRVM/par46rxX2j8UgJYsK9geoeGJUMREOMwVKdXccxT9bIfWj+URHi5G
YD3BMKB5FbhMN+JzVIERwCx69JnQa1N3y2qXahbrgCDl9eL68xxrbayDE474aD7J
ocAoj+3FpTD/Apmm+snC8z2cmN2rrMRkjiLG7LXj/pPbc34msOpgEPUzn4vE1iPu
r0RKiy3p0p5uiGMuTwIZ9FU/OuMU64KY5RhYkxbC5JOlQ/nrWMi+oK22b6kanRSd
ULcrFbreyIKVe/vbyfLSn0q1TYGFEKYHRMHmziTb6C8T0GQDkNFXLOkYtjA0xgsX
f/N8+cCDiuKo65+lvWJI9SUkwhXR9V0iRSDBAV4kQLyD6MyFJZ0joh/GmQGGMQ49
L4nRsJ+FXd6IBSR0Ee8d9DFYtNIvsajso7YAKm7N7MUNxQen6vLPeH8uts3VxTvO
jkLnagHCiaEZSmNP2C9fQPpsGurL5FE9R1D0+6ficLkw1omx+Gxn//DAZRL69jxy
I6ZgCGRsA3UlpyTPnFNwKxEfdj81zKUgmxn8V+qv9sjiCqiLFszeeTVnLUIKCYH0
wtAX4aJnbpogn7y2tQ8fPJrVA7Td3iRVSeS7wKniJ8zWijrzAUnD+ou1iOWl5E8/
bmWy9q0jPBmvhcPDqB3Y72R6FGq2M450x29V6QmekN+foAmtJxRl1N/6yuAouGMD
vGQ/CRMTCwqSoRJNKGRrah71vwxAkwp7srHolZ5or3Ogoyz5DoiwXS1fg39cKHRx
5FgF0L6hqAXcOu3vNZt1PmiOnQXOLYY9ZaG+HBxDjkF16cTBs7tIqLgfn5TRpHPA
XfP9fLb6eT/o+PpWRAabmRpwWYQktOd5R0sNCsCvB9OmnV4+trNyEUYnZrQ3weeW
kui2ASLB0LDJBTwQ3B+7xnj7F/J+cNa1+TGVyptc1IMyIFmg2/dmundK2yRJbasS
1eMSInxKg+VKZqvQxG9/S0XKQgMxCb4Y1AThbR57OfueaUMPk6wjM/h4ksijCXgx
+2kqEyj+USQztIv9vFBwkXubmgVxkD8v8YqGV/6b69edcbLD84XV0637mqxkocug
0i9QsKd1VwBbjwyYz+f1T5cCTiXIEQpZn4zulLhpnUKKvpxuTT+Z2/vOxGK7sMiV
kgODKXxZWkMqPkihVeCNniLEeGwotXfnoTVfSgRYpbqacm+nz1M/Hi75WVnSPmCI
LbeSafe7OgH1tDniyvm5zmhaE2CmMXFG6MOiRvwSQWyp42TPNkwJqOLV/z0561D1
K5SdU/C1o53s1EZ2IZ57joRwLHSRaWEhldjWsEvq/zz0VRDSz9L+Op8mHQ4WPIwW
t9mz5d+3ly2gwGcWS21X3un+ouIRWCZa/FxAWvgURPzLzNrhAktNWrDSi5QtfO56
kc/ftnPRUCMvDhet+i+ClQZn4LQxfnwCRezsXbheIN7ukwTD/o89hxxcQVkh3jUZ
EXgniBOEWtfg/94D/V9ALB4Go/d/YyRJaJ8BWtkaOU+1WQMU0UAzIf23/X3oR0Mj
b+38vffus0WYa0Lb4MOzzBDRqpwxYkV5Fu0/go7ycICzl2FOt3sjRob6q/zse9c4
QY1rcxeVYQbAK8XlBGQVvQXfE7QpwgAc3cr4okcAve7oQMPecG17uyr2H9wlQdNz
WkO46OWbRKoi+7uGBjwbKxIynY0yUpauC2uo6/KTJDMoWjktDbqPkRjtb3sdTnPA
bjoMx03xnkhEQhaySYRRxdkK1nbTNONygkmG5IWtACPoyTp+KVP9TaHdnJLo978L
4HvYAnE7mkwGCYrWzNvOsRLvGpC2hHn8kcHETaaHBLZDv64g1TJ2cDIFowWWHJNK
OFfzYB4R0QTPYP12CSlZRnd44RaTTFSJvrkNc3wzMYNg1XXf9iSP/HmctCDrRB5Y
qeBiUTO+UgH4XxYgjm84T7o0ug8Cf9+urTfQ3zdfI8qit9TsfXJgGosozca3uoc2
qVARIpX654mCTvaxL7++AfB7Cc0Y/U+iCqKk3NDZmtaRXPKHW/WHVvk1yb/aDMUO
nuct4gt7F0baSX8Uv3OC6ToDbzPLHWnc2uby9lZQLOpRAo611Cyg/4QnemfOwvGR
MEv+eWVX8VX18V+NxSRKuz/ZgFS5pgczcRrpp+R1kavfxe6YCn2HYdI4KLRVQB+a
h4+0VUzna/lxDZlX2HkZN5VVxlLI5TUMar0XudvncLKPt8qvppz/sXNVaJV+JqWn
NMbcmp2/3yvf/2RAzMhlXpSyzllYREJnWQEKx5tJZ1hDxicZ2Xr37DqKwAAcb1QF
rswQ3XzhNXeuaFoVwYSXjpS21HBWIZ8+KaR7YXoeUJW2uoZBQfq4jE35L0f9oU7Y
5T/xo3CSHNYX5X2Nz305ZYftQSb81Xd7j7pe/7ErFTh+vTpbCIks5ywlOv9X/25o
LJ2bIysBPdN3VaRaDsvymCpBvFQH85MlFf/2GB3kBEhTBeECHrAEnYwFAWNnTlIG
kmTudITiab9H4DIEmNj3+TQVN985sRauKtm+BFDr9T5IKz/2tVKjzgX4wYxYuTh5
FMe3525nC+So2FijdUe6h0vnPK/wtjfoK8wmA5ChPuz1ymRYElwnwl/ddWlACASh
wIFt3rwo0uWzHKmlMSqglom6LEimptiETNv4NCAPZCWLJh/wOkGMMmtCw9u2rmxm
nWMPKNwdpg/dejKr5q1FpOtAeNfRVqYhjWpdKbicuWkT7EyQycC9tX9IkU9jfsSv
Ygj3G5blUGTi/4R8pQPJ7iVg2QrqrlqoWmxZSVtAvETKdJX3732YBulSMvMvvedU
WTwtGzEeJPGKbYMMMTc6zlRFPXiwb+kCU6NBqqx1+lQKuA9VwcXSDIkSNObj9vtO
YzsesCqiksqUitWt4cUyDc1Pi7t+yQPXhavKhgbgMTHCfpemOUGHQRXXvCqKq6ux
baspFbmC/h7HmtDIJg7kl5WJJ2Rko/ZjTs6vTkQyJFiWig+maG7XkSfZP/eJtqhx
lmLJ8vAYse541QwoLDpZNo3d5dWLwoTc8sxkgJiuDoFrhWIdhV2zhywUaV9q+PSo
6DZVt7mLZgogFzDQ775Vc5ZqyZ6BGInc2pz9n8lDXNdm1+OBK4Cfg0ufeZf0b/mZ
5kzvBdLk+2chALiFLmkWIvhiuSEecokwUhR1EE0CfBHnZkJceH9sHClsU7bb7XwN
7u4dcEtEWMP1DnFpaVCGhW+Yyre4KAAdofzhVgmJk9QjvWeUraeA4ncMBoDQLpFM
KvhyapqkxaEn88uhebb005MJ1I7/uTouIPXcq/67k92SnBPfKukKdd4dIcFb7uNH
51K1lyjivnudlgym5kCQT/AYsRahH3gVaVNZgOH34al4tzPpTFQLbgswGHyjMGPC
ZFXbTwafkH7jq9ZUnfNF6UEl92Mrz6wpuzMddqhbPIN4cnHuuPCMbGSm0AQ7+TXy
AAF/sOqjnMWS5ZJ30Tc6nXilVwOURl1Fwb+cyT2wM9cp49fnB4/ggmFtT22Ob1J1
Y3J2R/krZlOJtKEBvBRJzIWvEDyqsDx6Ie/oe/TaevzUiwOlWhGDnw83AbKafJeQ
K6p0Zt7FpPQWAmP0xg3/A554lkgKLP39FvZw5/1YI+hATMvIULsm+4v5vBJM3TGY
SAZ5yK6pz3f8rYbsOUPxhh9tvkzN8bj7i/mb8hdPm3sPtNKLaKrJupi0dm3EO0uQ
/AS+n2hpch99vHnUfm6O3ltYOIE1/fs6z5sKg+PEznokYBjnFSNNjzRIJ2CEdDjH
ACihB2an2bNLxe+RLWdn5gYxjO5EvRRd8bIU1BquX3u9nvt8FQ/LW21v5xU7EeQk
APwt6RXhMwEmCwpG43jH+wbgCqlveHNJIHNfegrwgqcUCLpVKUZwj0f8/JhS/EZL
y9rEPaCxWxgFyXhfi2PASjZtoLs0twgG8jG8FPdPmC94M2XtYJE9EiIRpEQbzzLg
yCS8Wxc0QPaSDEGeu3pI0lnRVUSZExvNoXZHJBSJjYQ7basYtMdjFuOAStVtX/fX
JlGeGWJBNzXNKVkBTEBWJRJ2DDj0lwoLcvnNsL8t2OOC+xDfzkA2LJhM+mvPGeSF
wlGI7CdrM0ykY2jLTuwPjMAPYjItKnTmA21jvSETv04QWc+/ksQOZ4fhn1gqvaZD
siVTEmdAUgnWeDu51zDJIid61MIgdCWQyEbW6iMOzttQ+QYoFunjF3ewVb0XTeKP
7rqogo1e1n6uqrtxL/BDvhobWCLJRG4znmKaA3n0IJwyjA3AKFeKhxuNcZfnRf8n
FXzNIRJ0RGAXDuKhN3R73yOeM6T4RAPKtGYcb2+77NcC1eOiJGaEuuUVM844caJt
e3w7HfEMHe82Pxi740JPTgp60bfNEjRp8dxnLxTbEMfojci9ES9HILGzdwCIHHzI
BXIha4y3/ouEwhqOGLQEB58Q9gvbti/+VAhIAKJzqta68xwVLan5+RQ30JRnchiw
u52oWcEscb3tKQLulV99Hcn4E6vCdRwoyRxmxMlRmyDUWU5+v3oDl/J//i74XbIt
L1kwWBoSoQTEzWlGxMAvqhXh0IMuxjp3xmRbt8wyGYkA41DyuGsigAnUzmQ62UmA
Cgk5HXMs6WgUBRs8jNXEo4UXDGstUwXjrvZzBZqYgWJhkNaaSfE7Hpn4/8TkLSBC
hW5obQwffHaYgH1vm34LfegJ2Te/VcniC3YaG90e0p/RSfP7ajDmNgX+pw3LErtB
VsqInmGVNO9CPUAK+5SiDnZ54jRIq3g/brqCJ5N4RZlf+jb2fyNsrKKh0b5F3Ayl
58ixBgcor4rROmWCgvEqHc9WjQPxrLsdjYeOLOE4TUB2LHbvKA+nv1bIufG5Fup0
+WUALZmOXio1vEzQp/2se00FhtEP16qVcJYTAJ2BeEKBBPtQJv53oNrgZ2Puw5N4
q3UGkULXpWDijgPAFLXYzRNKq6h/2flHQdlqByzNQL287kYgnzc92WCOXED06dgx
W3EAkGu2wLhaHt8riYri58t0ITAYR39F056Hi/wJMil/86nFgQ3lzGBTk0tPJIpV
9cmlwGXklHTcn/BkH8uhDYd3Pw9TlBKuEWuTAqc3n9/RZg8w3Kei+AS4IoYgA/Vr
yJIBsnOSQdhNVXGzitys9Yh8k/YTM8AOy6tTsCiDmyI/xXn+Y2wx60hHO7hvPsPA
6U7T7+5L4Q9t9dyylyDWXTUeZ/BHHoGnhzJH/MrRFPjl9gq1UJl2yrpmpvk7PQ63
YH1HfI1PPZi5jpMSnO4WTWn6sLV4wTK452k3RB6aiDipQWgMrZd64QPUgjb309vz
ZmGIRjC6EEPeTrsV4R+YUkvoo1XadjiJJ9/5V23u3AiN2339+S020pFluNbLQqWK
abUIr7xpfFUMX5tLgZgxVC9L6rhZ2YE5dVqs1UM5/ihDSVuBn+iSt0oxIGTEx07a
w7dO1mqMMVFa5Bm/EqsZ7gCmphQ7xmuslw2HR5BB/qYHc9p6toEeDSwldQ7lffDC
kJ8kVtYynH+VX3jI73N1ChJWzY6IE7/Tn21ejP9N8f+O9pOaCwY5eJ/Lgdz36Rgo
LYoOmZE6gw1Z60lwhZbYqIIWXQ7YLmAW1F2HV6SWKCurD4e2XGynLX7641axFy5f
YfhayhO02alYHo6m4+DhykJVESEHOaVXlx38NUJGhcwBsgKfa0IkVGWdeICsZTwh
tVD7kg839xtJDihqlCw9KDw+SXRMYgWZEsbmw5j0rsvYFECmszxO6J+LuDpTAERY
VO5qA19JNgm+aIi7kR3jrvd9QMZsHNy9neuKi/M/ved1KV/kuCiUoxarEu4/trMc
rSaybf6ETq+MfmkQcqkQUUNNpemqsWqlYSLhYyKEBFXs5nvK5HixPxs2XdK6rflQ
AdF2p1LZFEc25r0JsaMl3Q6GEv7L+J2EX+aNwnSho2hWveDO8vlThg6PKI2yLFlo
LG4hkP+8g6fmhjvJghckOG3Xi5Egzu8YqTOYo2C8vmCa+RgnDbflH87FsdSnYHBl
bV5B+rAfrMDhkb6JxSuP6+Iy3Tltz3eoWEnsE63mfY3Hkx9/mvZ7NifLUo9dYJhX
U9udjMKn+FFdyabN1xtG+ojss7zK8XBZmkuvOuncZ+iC83ay58Drowwo/4ZqPjA5
vrVbWIBsrpboHTWj+/qXju1CDoXOOfsyMDSOZ588X+1Dn1x27VU6hTSNp+O46XYS
QAgXAfGmjiaagCvDZPdijpQ0+BisGqghuGt+eopqQWLGE5GYLL6vGhXbjiG2bPlw
Zros9YlVnzsAD/d4VFmC0545LLtX5XHdArzeHSP+LC4P98raFbLVAoBL2T7sNQK+
DR8blExQJ7zlSpkIbsB4b6m9B2tpuzwntot/eYTOwQm+CKZR161CaeOShOFUS/3b
XcgwdJLAhJ1Tw7bpCtmZ30Ijnr3168s1P9p3wM8MObsq9A5lL3nGOF4fcDhAup7j
TdwM+SZGeaFBkx2D3Bh56Y9VfVkozqQNHutqikEF/g1u4MGamHQ/GMd+9oEwiLuB
O4EHTZA1m4T5nwYXYP6eZlvygCG8y/8jo8HPaLRQ3maywA5Jgr4oFBqn6hDzUBVU
TuZK4NThRp+CAvrXUw6T8ijkOhfJheZM1C/+7Ks7RUgyCjC4c8YcV0Qr3612iR3W
vt4DWLFUEBtXbpd/UQyk4upGIr1+I4L6akw8d+TsevxMFffjpIMymyFCUzARK3f5
DawKHX4Re6vJ0EkaJEa9xbOmY9s32gAbejKAoa5281So36UY3XnRD7Xv36FXLz9T
JvsUqVbkrR+yZlhefuqSV0jQMvKnEYgjAb7wDG6YZwzhOaUyJuNPVfeQIXaOO5RN
vCQyaoqqfVNw6g4UZqyw4Yuii5nbfn3znSWZ69YlYw0ASZ/fU/39XxqRRGmXsU9U
uShaKVH/0l0SBch65Gvi8k3Fba8H63AoPyzCN6WFp16mKxxte/JL4eENzyrTgK0Y
4UfoQn1zOgz2ny0ThNVWngzeQmeZmC4BtKU4Nw3VMWO84VcK6S7mRVVLSfsJdSCO
MZLx7Y80SBdbjkKCEGXsBMBORyJeRtrl5IDTcFqOyP8lCOVaNz7R5j2aSPS+DrSa
6d9UJK9CirenhrqhN8HFQXnNgDTQa38sQt9CMk+YItlNz3OlxYiQrMShgmnqZSOE
+TO7dc+ljQN41KYh1ORhk355ITYL+nsQaaPzxa7KlVRmNlckDRmXycNRMfrRfZtT
GOxyHN408XNvOeFtlotaq9Wlg91P+MuisGJSDDk9A3GtmOkp63uGL2Wi28OvVCHt
MtlH4ruTB8YLfmsqXrREN+CqSMXKCyrD7UD0EGOAAC1bBp7M5yxU1PPsG0CugYHp
syee/12Aynjt/aMpNh9mvMUaQeSXqD9j4AztwO+MeOF43XLqlvLt26bMLVceADAP
kl2lEmN1AWFKhHMS6k9SwzZ14bl7/dYo7p+LNAjVlTucgesldqwkEJCqRz8/jSwz
/Bmy8hvSD7KoDNfyY1EVsSim6Ax4CO0C5HBUO1yETb0NdhFddXXVeIPtxaw0W3og
vVW00oz4BQKZOBRA36ZI7bZgfaMEQndgUCereA1brUqxjYqngpzDT6VqwHqZfCiK
0rzmXiUXxSS5AgxE8akfyCb96PJ6u1POggrplgGOqQOfe/VrBK8FnY2H2EjXcmDD
WX5NH5LPXoqYEqfo1QiPHdwuZfeiNhj6xC/rYOKPHIIE0NX0MFWgxzgWOEHnP/qU
QCvlV4eBnKSejFBocBTgTzem8prUxluL3yDcg3A2dsmC6/1X0HDzwG1BqnoLFinj
V5MSA0przG+v1gmIm1AKbK3X/0q5d+bywv1lsXQI79XHBpwCcND2PpyCAzls5p7i
/y5cEDM/F2xg5M5he6nB8uJPxT6MKsQQJQNNoDtA7sC3bfWf64pM4SerI5wbx1Oh
/leh3jEnTuQBs5w00lqmUJA9ytWExBVLfmEpG2L7F7T3HXixm7g6hiYwxp4C5NmO
CUwo18aL74X4u0OeqajfutKuLtqY4H9MLjMew9fO4yAD0zA+1n37vUXTV9azsPhA
LRcLjYgSuDt+C9XcB/36FZFS+/N8GZuCAE/TtjsWvi+6RzJ1mxXBj4ScWY7a+Agt
YZawwOW7FZBUnrPNrf4ERflTMUeXSTXTYRPtRPrxk6q19PlgqR87EjIuWjwkeHNy
QCObK6g6jpjG1rUYmU3xNQ7gyqxDngiIf1u2sJlGv9AJL1RkqOaIz9pd3FfSBFUH
8giNxgjDKB/KXpbCKrSjMSbgn4UqVOWElLSilsFZv7e19rdJkvFB7ifTYSlGFSWO
jvMGkInO8nlwmPTlrig/0wOx4+/nE6IvDB7VnXjPpbDu1RMJesnoqlYrQvVYLgsI
IJASyZej312Wz7w8gEaS2lP/WBmpcoGt7iMNbYNBC6o/Hf+vsRs84Mr7oKfzmnD7
t7+4I1UIX3GyjSqpH3fehe+yIdJmCtC7htdMJrXYGUP3zfOLJjDHXKw2gZcliArb
fOZ+VpCmlYEgAc8pClS6M54ccbkMpPweTc0/+FvB9/ss85yp5phYnD2GzUc3oLZs
bGb8iTgU8tanRxASgUojwPdHHCf5KXXgH+N4jSIEPaOXVnGRiYkpNp+jiCxb28ZD
jwwASZAyOhFz2RJgjBGv44QiN+xUf3J9z+t9SODCxQb6mbMEYAazSvw6nfBewKI/
kcLxVexqjHYoX7LRjE9dZRHLTEsVOeJKZyEfqFQu+uPfoOpcQIFOoYh87bMKhipE
e27AES8RbOVXw4B9pGTzGSTGbIyyfj4ljWOO3wB0kMjTlmg/IWEfPRqwvx8yCeJn
BuBF9ftK0fbl4fSOyWQKxFLSreHfm5QJEaNndNtP97OR3V63VBcPl0JANpCDNiqd
WdAKgTNEuqoqxSfn6yKO0t87RN8Xj69eV4SM8UEbyVdxVPVE4mKCUIDR5Ggcd1NY
3RZjKDOc/aSUy8X8IABLw0OX8gcO7z6kykNQVBTORunOZjym+99xDRaEzasN9dl6
o6kvejpfcAYm96a5hmFnYok8ZeAWMHCBhdhkCBPzoEtwpDXT2/1kkziqp/XgxqBy
6IQAGJNN36/0I3t/IQ9grb/AnyZHoP/KfJDOJ1J+dNjlklIOn5lo5YeONaSZuBnP
88xq5wLH34pkUhTtZg2cBsXkB6F+LbMZnmP4WxH+dGBFcDPAK25H8RlZJ/oSLapo
Z7wcBrwU6euTv74pSR47OEZbI4fDnSy9syD/oGyHaGsJB3SHXUTYu68kJR0gh3F/
wPU83mmxBS04gxfxeK7sVZTr+6aJ4A+fhJCei0bUhzqdJle4f7Yfu/ymWgxgYsaG
ILGbT3cfl6pWHmq1QLYQlaDE9ZO8Zo+R2DkMcldG5j2mAfm2YLlns7kIHbpr5QI4
EGYfxQ2EWrQvHCB35Wn/DWb7ya65X0iAIZuZ38RVuE2AHfUAGeQ/pSm8Wdjp/Gl6
y5qd82D1SBLyZFU+vflPb4MQjY4/oE/cQsVNrfzQI+RS47vDyfpxkqN7uh0u6JGu
DstuuBuGCEjCTHFpXusxyVf3BeBs2PDGiXiF8JLFwQlyDJbd+ezESpyiOUJgKPU7
k+r/d/Q+LaoUAries9WZOcWGT97ZRWZ99wZ9tCIS86fwPudQvw6euVkp0SybDMBj
BOFOIf0DNx1Km3/j5xHmxfd8U77bjM5sfK1/151mjhn9yE3hyC0sqIFfv7hDNlVO
OtlbbeJ7EjatNZQO4ge4I+Wg2iNjFHwrL93xbzFD/p8ZvUgVvU6MkrYi/ytIg7up
0GGxdqMetPsk9tc+dq+ArUCbp4LpY9rNLxl6AWgs85nAWdHrzO6zskysK7NMb7wK
GQNcyz0dOhwswrIlRsn2FbzOlNrWtxguugIRDDq5txU8dTHXkruSClpN4sIUuZjt
GJZcwAcpmO4vRRYi3sRM3iZ8UVfCRHXJANwhHQE1Fze4Y72BxLPNEVGJrO3QwI4Q
B4k6Ic/DfuCGxtgNRxTpTKGr2GBvvS/uiekF3ztWdreJJ6ey9r32c4ELr25nLjRo
z/NmtKorrK37vitPdZZLfCjnNpKxywxQMpvZz4zBB0VqqOiNKqpEMTcumGoEPFJQ
lWYRSDqMkpq+UYYywC3u7VKH74LcB5llvczUthmp54n4AEZb3vnhDAbetTEcw27Z
yWKnt1NuD6e7V3e8nZ54NvoaltujSHGW4lq6oDhbU2B1ogMahRneZdgmHmep4z9d
yoML6yMCa1y8Zhu2+fa5gqZaqmN06DXiPAYLQMU8T0lEsCJ6qMswqmypX+0n1Sc/
vy8TfiVflm0mMMcQx2aw4z7V38w5tB9UiGxdef5QCADjV1B4vyw03vyhV026j0hL
GS9caPKiXaTmgdU5au9xlAu1fNl8TSr7Y4wOBlRb8GXiIhY/I+hbM5FrewEN+Y8V
n83AoJxiRbCa9sVffLMysOedsviAkOanNKg+dxgVYaf/kBi+5MwbJQVANIaDZpI8
YTyx21DrWO1zr0oQNhY0fZmhI/NTdxuYu5RXehOHL0cUAzIDLiAEMCkiJXmTKhJA
h6bA0s9AwGEfznQXve8luy5yg9Ark5jyNoB5DLVWzLJJ6tVjT11KV2G2pZJbr7P6
TJrtwYuwDSRK3YmbSQAy57AvaLzxjbdvyJjJRQmLdhTrNW1Ti9DHcQCknTKhy9ws
pDz2BtBfZD0K589Z+bJ5pRnxAtKL6XvNcCmEx4dD9ks7YkXn5UkA8UgRmcS83tiK
gkeE2MTg7iWEtTK5WOcldpOB79G7v1XcPqSOyRBr2OCD9vkNxMslDKktNShRMSQP
m5bv4hGry0m2JZTIlwVmXLhyU1HoyOPDhac2CuNFXpfj5ZeZ1vjcVFtejDdckSfk
AUhuQ649GHsIZB9KngBtmvgo6SAkhzWr5a5NAnVeF8qc04Pn8YwYN1QrBfkwYSp2
sY7iJdkimZ4D5z9aP2wcT/fAX83K1Nzr1u2xFUwUr6CHPIrX6ck4zctPCdW49bOS
WlzsCI4anqXjBSROrAtMSVmzW99CQy7vttvSObzgBfrv4qTETkfbQjDvU8nU3zOk
rEeAMS+vhE4h7SU14CJNML6BKgd8YsSVaudmA51W0SG6epl4sn+Vwjhd1MSbU7Oj
TXE3Qdhfu1sdncUwAREyl7IwYUGVDs/HqyxW4jr7Qe6/G6ZAD9sNIaVlDxJrDL5A
BJcYQzm74wAdxyLgt1lBHYNVZFhnzUsrrWySYNCwDJTSIOthIWH3zw1g510pHqWI
CUHwNYgg4Uv0L2eydPvnMkDmBG2m+wpcElsMxueQhOcLtT9cadeCnk6SdLYyHOJp
GYmcnh70WnxFmanKsiqg+uINlGglKeQnKmmWHg5iG1IVCCSE8+4ZgbhTOajw/5vr
xhfFhnwn/BfbKbAilBx6hFcLlBwfptXDoVdXhmQhBJnLq+fwif2eT51sBeX2aOtM
0NysUeKFesHpj6Dtvc0Txmzq/qxbimPnr1yKV16Ko1YhTaAIaKa1EtuDyTOZGPUG
ETz1EsQO4xcpebJZWANJADCZydbSyFCrZd71XMplfy5Hc/2iA+vFV0m4TYFrcAOm
R7R0gArEHnWhz0aSESJtkJDGjnrl078nxaa1RvJlnWrjUsJx0AhmF+lwpQjQFzyL
uHfOUSPhtVgX2UW4s9wZmRhUie+XXSQ5bhbhKAf/waMqbZLUsMbpxHegiqMZV4wD
czLkknPbqybq3ouklScliUG/Ofi2hWJkohN33+vcx5Py8OPXfiKeqNdxTHwCjic5
lrRW/8BbgZvyLGUVrZvwn6BzZu/252kiHc+nKBos0zDteTkeUjE4oxeK1yNr50ij
WHbWJCikiUwgAOZzkG9o4izrVv3jwr97l7JPq3eMIoRkYzzLJmVLTSdZjQ8aKmc2
VhKhrTucBQNUJeWx24rNo6LXieN4R4rjduSEIGGDj9xZkxiOeQFUsTQqaVqXVHWt
HR/54U2o2dpjqhpI/BbWiDpsC9hlWbKzrnLmGD/g98w1dsDGJoUAVqbBdYcvxtfR
8ptmoXwVwvdvm/ucd3XfNtiYXAmmOKn2WeRxFQtn2R2ZJ3vN/cVlE8botXiV3AKy
amRdZtk1/+F1q6apaaCZubXwKmWk6onwTdOYe9zE7ugRDnOXsKZNStvCOho8bVkd
Kr7rSXrxaLX4NTezXqEcNxnOl98OfZujktlpDakWpQDsgAkc3ypbnugx7UgVPRz5
nhHDltJogv7Fy6qJgIUZC7EN2BRwYT7DyZyd+Av1bPghESJCArNpl6YDEOdVtzgd
kvGh4y6PxoR7lY9HvNPxJ37jRDLMStI0Gjnw6GmtkFdCOAh2j5qYs5EaDNqJ4+Z3
MNbcKvZoJXKzJFB42QMrJwIxDyuJNTNvz2Ppxo5RwH0j2u+LQqb2AHZ/KLKhdYyh
Uk6W0O41BDUxcBXG/9hKSgXyrCXTslmwkA+1yR6k61IPo7n8NBj63Ylz3b/5Co06
ztbtkGh7f+beBnCILQEvZEIwvxxjrh1/Pdbe3sKBIRxszH08484MnDQxDSCf/j2w
4aEPUwaXkYqsiznb4nQ9pJnNEDP2WSA4JszcjuuAq4djIFLtV7PK67hBsLJiX1sj
VRzvT4ovCywvrf8OAhk8LoPRjLW/HiZuOSy/Ou0I6NgL1geJ5kv46hVT1Sjn6mZQ
ygIUlfUBYf0mHsCrYm6jyJNNv4NkaRgX6ZUCbyl2GcLdlMJQWVA4/0ARQoyXAdu7
3neLYsv/hXhMl7eJT7tlgH4/okqiAm+K0J6aGS55Pt0tfhZ59GQY6Yqb8z0XW0y8
f+x2pRww9iBTa2gp2u0Vht92eZ7KYgVw8zh0ZcXEMHd0R7KqxCN6SkqqNgN4Taf+
+XqIqIPiQ1upkGMrui2XrD2I11v6aVqWFgLyIk/QYfDm9D5Kr0ed1wUDKS0/gWD1
0Wrk+qjDq2P54Yb2SOOEde051jHnsjV0BWA044UYkbA89r07/t9qIOv4V+6MHSy9
+iNN9SRiSvwkaofb0/fD2jSNNfl2EAL9PonZ0qwj0ZThIE+2bwtlpXUaFbOzDUwY
gJQuTNsYJ92G5ERuC5CWsK5RGGOGUOc14uko7jrsVyZYr1+oZ5wnpaGAq0OMNTkY
oHA+YpbXkZYxAxRnlBK9HsRdHSb3SaRl5t5C7q7zeEKbN26v/yRHKCrLWlVgoINn
koo1c4fN2wGpjKH3eAvB9pU6vTMkqvJ3LYAH1cLNc6ZUjmvEmlDZ/kXs3hi94BdI
VDgM3P87yhmBytZNzwE3dDXEhODHThRyGClnZW5wSDvLU8OZT4PNXt2Z/r0kbIKn
R/q0nX77yWJCkfKHRoGuOVThs6mek+WCehnN9dGkmOO0EScmPkQw0ONhMUJPSOVf
N/JzLLfUHJnWEPKfGc25X7pU10S8jr6PVmXMo8LPORoxWE1N/KGrPzeSoIDUse92
5e0cXpa1JYwn9nmT2EpIoJK7bHuAgl8e0NOXNWht/x+lOo5aPKr+S5/laWjz/4G4
EA7jqgoE0BoJLBZDCinK2Q2bQQSmML25mBZ4HMXO06zo8pfTKgKBLE8Affu1H1uG
cJonoT7eLisyanN+pY9OEHSayI17C8YGWgKDotO7XuMtpoX4YFdUNfeGuKAo84Ud
24ZLNoNIVfRWVXgHNUWMe8JPEUkdhKz1cnsSwShT63mlyaJR8GzgUz3jF0K8X5NH
HsibXO+gltZNaIM2uJbXNk5ppDq2eYBHSg9LnFshwsddPo+tLpNYfjIC3Vm0SAFf
4pErsY2TGHLOqejqdRpw3TJgnFIhTXbC6ieCSa3cM8Vqs2kYlAFBgdyGEg+QbM8h
E6toe6uRoBXFSukrZywW/Usab1WJ0ea9hboAaRTigdutaxWKglKp1qwVcPbB7QAk
xQshd6fMggQoPKSx6RB2b1sDpj9F2orEAkzIRSirWQpSaCQewnPK3nRvV6livrIV
4z11rrPUURzQ0MJhd6A8KfVfZxOmwGZ2KiHsS2dns1gktRJxejf5Ne4ssJCilcII
JJp9nQ07/ooiv54c5u9JP3A4zsfLtA5ERrme0G/VQ6C20Bx6yVKvnl16oypOH0P/
mwm7SNBpygoAYaqPkx3g+MM8yDQEmVocf9dFLtnwjtDGq8/g9UMU9r8zJbUv7HZG
q4ZHVvQPTjdcY87vJKHpArMumquRIAD5PmrmT4OxYRMBVMS43/cQfSfcNY9q6KOg
nOPmf1deuA2NV75CeTPCriP0B1tXqSyX6LxFTxU73QVvSHdjmOWH9Y3TCcoMJMi/
aGywr1xeBWUSeof4pNIXVhhYO0kM8wYzGhXqTs/XCL73HymxlyGgQVPqmN4efaeQ
Y/s16bO16YzHWDCx6SIF90e0RFuiqb++EsfHbsdNftMoIocqA3EUWLpLd9ijokAF
w69qpVZoHVRfbQbf68Sx+u+NDjPYZIJ6Z79BZomtqfWY6h757LCl1dgeRGJOoi0D
w/jWkxQirHPFoIkv8z83Uc+HPpnvHBPiZ0qkAGe26E0xZJGmqxIWzvj7tiAvto7x
Tcb3ZoNypZ7gnHcWqq6DNO08K5NW/rmKWiIWMiDrWnvSGwCNUZgm3UuFHExPD7Cq
YJeSS4Q2AP3aJYqkH2eigxViukb4EcoRFYvHAkdj6w76HsjZljmrolKqqHpf6SVc
NQqW1mcmc/OyC8Le/x1fY9/vQFUkdvmYS2v3W9yz8coPy59O5TX+XKmaiy3TVhaF
ekqNKE95r2PaAxj5iuTHGttkv4FD3fi6ujSze3TW+bmSnH37MblAanBj+U5MCQSA
sHQuBZN/bmavjyzg34xdtFGqsn6EwQRD8qqnx47Y2489YHxyucVmbFrarmD3svnY
QFYcPz1qjIet0fhemyKrosDiUNpV+oygxCACE39r51WxkwraGXmJRw4aBMb+wWjz
psSmL+msP5D1BM80/6xduM9pgK9f3MyCbPF2WV9wv9cq+k/dAsm7wiWbJPkFOrH6
5QVMbmQDxRzmRTliEE3ENQNtU/1fZ5iwFYN/PQm1Prq7QrFZanrrZCQ44MBJWav+
XHWv79r924apsYSXTgahOdYnuvHD2Gisj0Uvuh1MoADJK+b+IU5HBPM9DBUnArKm
7qFVxkY8eIRIa3TZgNAlDIod3DLNMrj2Plh1ih61Rn6O2vImywMty/x9IGmdwoL3
6gSUf78vPU8TRE2bZcXjE2p8IoARKJzkTHZ9exdq3rqbHU+7LCPQfio4DNcwUjEo
1KcTDvtvGOatwjy69QTzrzfpuPEqUqHvhYlHyTh7tx2lrcqwdmjAELDj5+ZQKdzc
KOTkC5wuQXzWbwslnndbSeYHmlCY/cjwWWel7fzS4xb2CP1ARmQIzly/V4GQ/FGc
kPLVXrRG98pnxQHmNu6g5K0hsy8qHyamNkhr6hZb6JBQucWFibN3+rGQ/fTyrx2z
yFQbNAO3DF9niltk7yoa7imik1OoWnbLNvyf8i64HmLyGxpLJAtRl7XNdsqiaJWs
fWgRgop5S5bykxrRnbvV3bs+Qqr+9Z+erV02S/tsP5yYmLejy3LugVnBaJ70fFrw
jk/1o7Y6oWGoNkzqMKX/6elJRHIvACtu4b0CERnDuN3rKShPpnePpsAIW6a+Dbil
Ef0o2UreV9PGGSoUg2quS+TeSqRivEbFwNNr4xszyu+XVI8mwOx8iwJdQ0M+31wY
BCbUvH0hv1Bf/J4CMZxyKWJO1yAVq7LJUH9eV9q1tBuKLBADTSB5QDPBuCQ9dyzl
hASLrWQlh+BO40aDuU+OTx+GinHTjVMa69I3SHcm4EIxKjY++L7oy74/W2vBppl9
mOH+62OfJlDEJcQIGg+sk1NM+q3EwRAQy0T8k/b6+X88hQ/UYgG89eFQql8ED7C9
9icCX4/SMz3HK3hy3kRcDcdBsDrlHkY4doXw3gK52D2fgzLXbZJB1EJQMUbx5Ljy
Icq1CKQMbrKmIr5Oe8SFBBqU2aBJ/9EeEkNNeeV/O1mmMLMRX7ybROPUrIfnPM83
CvcLW4NANS+tAv58IpR8n1gdhO67MhIhs6xR/e/9iAl0YnrY8WH9T2INLwJTmJ09
5IVzOG74leujQkN4O2UTriXleR6XmhyjKN0jnRmImSKioaftDM2hvElZO2RaBvxO
1cwL+AP9u6lrpyFNHzKEUUJDUewPkmz07xC/ElgkuiDwcKhXGw/lqnIkdZhhO5Z4
CkwAawbWjoZV1Znhx8f6KuwTJV+yy0LdhJZIhTGWzr1qhHh7hMEXu2wHymOz/5QX
R8nuXDFnCsoABcrihxN75lwY70EtjTD5F8cmHaUxlcdnw5ELJk7ddrToK4HiTKTd
utnilx1RJA/8clFikkasPXF7bcRHKJHRoFkfHzMwHfVQBrUq80hFZ/MHW663gphw
Kq+AgLyY+toDFjCOyqAtwDvLgz47FzMGir/LO4QVPTo8jeIqxq7OhFfa7kV9lZqL
eED+Ymsuroo3nMFAA1VY7o+8vos1T2eHHykWuLc1wB+pV1FNBVUWYrgnDx0wjK63
7tb/3NuWiePgnhFIS9xwNEJoGcWENfjnWiDzohIeJ7CDfGtms9bivmFI8BKCEyQA
s5mCPkJIAmjqrTW7uDcVovVkgXgglX3Y/JfukiR4nY7OVNEJB7H4KT9nDc9J7cF6
+Q3AoY174dBDFqu91dyIY8tSZoxdbZQf4xmbJq/y75TnMZiFSxiixx91vUBZFSTl
M23ifl5ps4gqG4BxT2wVTMVxFOx4UVUf9q/QdQWgy4/fkALcU85RGMcbsNTaft4A
j07xcIhxhO6KJO+oNsQNbL8gWEq6kxHgWT7Sc82JEPAx3sJfLo/e2scbRbjiamn8
79R0Pc4gVqpHT8tI7hkQU9rgMXO5ve92gIpOLR09cBUkkFHDNHNKvDemYV4tlwnt
9673o2s84d+BfbofmpXaZhxvMVjRTn4xYwYy5CxAxB0TY5VbfjoviIJHGN9Oa7iB
luolCQouBVin5Gc2kom2UdNH9s1L0EAQ5cFFbdxytvyZwd4Mxk/+6TX8MWQ2UTXf
YCOsakvCG7yY/djDPb44b2lOKUDoQ5aYhSbHq7aAPibPTPSbjMx6RWbnR5jgxZHU
y9L+PsE779nx9ilQKADpvV3OjhtvJhc/aEgjrtk7MQKqCexZvlDQJ8RO+2gZapIu
ZHiG+wLm3Ll1uHdNurRCXpnkuw0UVScdvtMXLP5CsQgP2mCdNqiQnTACYciJTiLc
lHvmfbu2tDuFsLNLzz/DBISXMI3eZLsf0pb0VizYoWAmVmExb6TpQmub5HadNeqe
NM3NeTDzhhEbTGLqzsCTjuNbpX4Y4S/8I0Ab775PE6aPp1iMKyRpepDhK4fS3/+w
cPZzLzocbEVnDXVMYTNTw9/+tuRLllbzQ0TxMgDYFjq5oqrB+xMIYTevuIEIu58c
yuUOrL/U16zM2iyt0wWpp6bxgsEBpMVveXUIek/K4V0c3DYZV5/UDs9flsmDYsnL
Ej8SCpJNHhv9JoRbsEaL0J47DtZCILMwlhlUB/sXTbY+IL+C9gSUJoG9a6My3T4l
MakSwikN5A1Lp0/OS9CE+pKA+10yAV0QqYC5l4wsT+fkRUdSUFmWGyZjOinVvcWQ
2tyHFbOnJTGk+hfS0MJbteQMWdKLO60V3zwggSSQqgFs1XmjYZHvlwadeKid+qlQ
0aXAqUwjd5TDvwf/UMZPdNChsbfHQGNbuqRlYcu7+GChEQ1KQFFkWCW/Xpc6GMhD
9in213SG33RYTTlvHmhFtHUp28GuMWtfXxSa8KSvg9xDwpCRPY9S1NTtFW/oBD4q
yL2D2vNTjz7lWbGwYC2mJ0uF0AL2TtHwxKteqRmTUNzrF0cG6xoQWHoDJyCNL4lR
HJevI7YC6oPC6khDTT3vXt0MG7zcQu3GoEBOG7AXqWvUchKayK3DvdrbGpJnTOLH
AIUCIHZqbw67cixUm/qUIpWFyaOb0dHei7rXDr3n43ghgdkhOCmOgPtV2XpIikZk
5OgnCAWgesXLngVxjJanlZcOimsCsi8sTcLcXzSjrBtUHMYcQnikkTPsOlL5rOKS
s+O00xVnr5vguxllRJl7fpRr4PDTGQukmBV8hiv8S496+MTZ5LA0CXSWbgf83c9a
JHCrX/ENYvWPCrYGJpWxWKcr/B4pv8SHpx4gObLCQat0Ol+kJRTJ2hwK0wN9or96
O31VZ6MLVaxekQ98vFAADtlSrQpXjQSzVZpMfbAwEL2WlZ4fVgiaTy+wHJzpEYOm
czUFkQWM+iXM6rvfJ9d1KW1moUkzVxdX2biVGARfkH8gLzGuWUZdzdYmUicAqxgm
w4YvvJN2xhVR2ME1dLdYP0QvexQU0PW92jp+cPgv9LBjP2b5M2JKrAZCfYBFwanA
2IJz2yPtpPYCJNRxcyC6mLayFpNjaw7cK5igIdhFn5nR03PlbtBWqHyvDrkF0wWQ
nk/awfjR+s4cgNSH4veTFb0Ck0O+ubMfWA4TK3TE/CipodwDOVFISJYK+pqcgzU1
zbd6zh3T7rDu5j9ojkH4og58urIKjGVUx0paybVQsF/uP7NGLHfbtDUw7YHgECDS
b5VQPKIUrNRRefdoByJReYJCAcZOW8EXxfQRLYOPCJ9vQMCe9vPYEF23Z9nRy5AW
En5Z5Nz7Cy3U6gKc10y0mLQIdKqw41rry+9yk6d4Sm2FbLvIhaO50RTZVBKHnujP
7W+05TTk2TzoK7cFiztuIfZbJenkKpAZqGfbK7cmAlV0OUrMVBdFyK+zjbXrWwoZ
2ErltJqmg8XJg401XatOj6tvoRQ41e6OpcLNBOkq3yarw8jAQz83gItNTJTvaE6T
92nX54cI/GL0zE9BKZUEfbTfsXrIDQStwzSIxdHY63g9HSMW4eOptSVrm3c7j8X/
m8qJz0G/uysNX/DX8/qTkabdzG1rTRrf/zDdqsyum52IsBoGtmoXSPFOtHz9m/EW
wyEt1r0+aWEiN3RHJjVll3BSA7Ei6FJ4rpWHq/nOH8z1E/ZWpZ3K6x5pHfsM/MDT
1VJEQrt8Eh7QE+ojkqZxKFcrG/4po+PTUcyyDE0oPYeWziyvvn7OjFoPjky5E2C/
xD2slcfKaxvpRZBHo8H7LLPjvbrC8l4owOWyafOGIjKKy0Ti5W0N1vyFcROA76RZ
efv/JJCHNbgQblHbxGaQWxfKpZ0oQ4Au2VjhChN2RlgdlTkUvv90QiXfc8NaJEhB
OBSbEkTOFd894I2ZXPVogo4ACcdddhTGvzLv1kGTRZCmW5mbA/bEm7xzGNnIqVtM
l5MgFl49V/frHjluTPKouzBqtkrCZ3Br1bUci0WpN70++/Styqro24pLWtl0qwcs
g/uFzNhoIgcIScV4+P8qkbA6XnIBKdV4exscI3Yp2hYjPDYdi52XUYZGchoeS74A
ylKwYLhoDLAyies0KpIYnXOJOXIduhwPZM+4FNI1zwD3KKdX5EGSaIQWYit/Go75
TK16CPY98F7JN8pWDuaJ4OCScruNmaJfKnKH9s9Zrt/5xz4Q4ZFx9KiYvJeZU0Pg
esbCVdURrD9m75ZLCFQz8bITiUBWx9BTRPDBXGWnXxWeaFFxxJxAurqitfabFVRP
2tO7MXA+8zmPV8pr0zxFmEFTZkXJKxSHluw8lAbszRqIM7gsbGfd6lUdLFfziC9P
PRpkgGm89yh5RS2XG+Wy0Y+IIfase95NfeBNvTZRs8mQxI8ipNIqiu/SmDT/cuXs
7XZgg3hsa1G/hOOGkaUUumSAylxcbTjPP26Hh+6FC3qzWurkYtksIze7AT4Wd311
8gu/QMlNzVAefGCiBfOHWgrZA+ap3sgONDvuMzLVU+uxQZCr7jIIm4aQ913VqG5C
ajsiz8xxzr5ZwoOd7gN/O0ppyG44/6EJr4DzyOPKgdwBmAiPb9CBfn7jKImTN8W+
V7n09FGDs9vaPq1jSexRs1tOFY8QRlB27ps5g545zoEfzxntucanKqn/h+2Ouom4
9bb/nESmwOYEYWKKaNBaEgJL2YgKntMh/B0iM6XAAC5WfkPLPWx+M+I0HY5zY3PB
V+BwfRgwae/ztLFhyn2j8bv+4l6UzlOs4ckfQVkxf++j74xDpav0Xi2n3wa97nsc
uExfRAnqaFgp7nL31pMi5qZ+iW8bsgL0fVt1mxXLeBG8O6X4TQU98tUwtHI6WAH5
SCO4ljpNZF46jTG28QvJkPuCV5LFnkxpsCNU/gbZ+Emv/jG7qjfEOradzba88H6U
GBNTp/xfm1uLHxLoFSPcukOyGwVIQWDfVAYmp9gJ1a7bIDz03d5P7ZkU+H7/c0lV
edkF93voitwQ3vABhaHBZGPhgYZGkFHHvdJ1/nXFaHSuIBpV4mcRhZP6l3oi0UnG
RjPn2/WxR2XgRAHG+0YPi0iGfwtuuZK+IVbKJCWNqCdseYT8L8QNeUtWLnTe8kYT
43fhQSEg0JHoPQKc+Ne+py9jJEv6LpAqTCoXCcF7tKYJvYHlKxKtI4QC5imJlnjK
GXAXeCgRe5a4IXDzH9jWyiWRFoz5t5guU3aBbNbyqm6TItqguR/pLyOkKmBfAEBl
aGBMwABc6gSDK7ARruzqeU3Ae4scGl4etrtqQ6AWHlcr0di+My5S+BGfh6azTmgt
9u7zN1TQTUhv+I2wE1F5AcMEAsdSNHdbXLaZ+hiI50PFtKIRzTgG0cJNQVggf4Tb
vdeIN/3+D0urSjuuvKy13XFzjTJEEMMZ+R14mLvYS3BQyKZgomdOzfqQ0pvgtKR7
8i/7A7khnotH1BFk/jMLwodaGG+7LbvdNeTaobIRBYjjsFfw6jyWq6xikDF4SIJ4
Vf2NJWBDii8ia25yz0Ca5DD3Wjsc6OogufmqlO4ZZyQ7IvufCCLa9QCHQOaiDWwa
wEt4GxC5no10Kiv4fx8xrBCCW9U4loovFV9srJHHSwCGv7nYBzeNUzzpfpgX2R0k
JuhUpfIvPiNjWvXG5evhoWUswmp1RQTJOKtTmnY/J40WuMgYaH57EIl+L1ciU2Pw
jqOZcZMDAmcONDe24bh2C9rqAPkVCEAadBLtiUcYC8j75ljIiD69JcbfRPEklEfV
L6wXwsk6zXYYOpYkrv1Uz3Q/2G+uTgNsYfqtMMF+7oqJwJ78eLyTBmoQwhRW1i+Q
f14C5133q0aAqyY6zUa3ul8arLKLOcUyxV1Hdaudr4zWKB1CVy12dk1Oq6B3zcUu
Yiipm2NOYxi428qn5aubk8hYbmh23g/l10UTLoQ1G7FmaCIWsedYtACM6weL+YPd
OnMCGRBSgTwJsI7yqwVa5It4yPLXnusD0Fs+QKEkOoUGyrOznrCqRfBP10dzjLfJ
qgRPw0qfopX+Nhj1IkbuSCBhsm4MeNMOQVEn02/dfjEtPA6U+HoerSSpmIRhhuue
5gf1YCJxLoa0ZeeOWkrVou6AtqIhNuZ//sd7DffrCBoM8Z6LKl9nduZHOIrziL9q
LZNKTYKvP0F4XcNwha2aCsA2iCZT+t07GDnBkQDjKSvYJaI2O0OCrvom85Euc4Uh
ixkwVYEkRMPJ9sPHv9x/9XSVct/4m9OCuLmLkVD6wkXBzGyoudgB9RcajKD7Z22I
MWxgjTBBHz1BL7iepybIVzJU7+XscvV92VGcqRH89FzWwFnD+dVwFfZfuSgRJN7r
RvClELlI4Nkj2md9M5GlqWpcw4iJ1CMmm/CMSz85pB7hfhcx9oqVb+b6VTXDCi64
Y/JAmerlT7OMlCuY1n9oIAXNrkdX+Z6DthX3Pqk4VRIbwsz7WYEBbdPqdYv5D2U7
z2YzNpSHUTbZrHhQUtuodsGJuInRz/kO2P31wjSHtq+6Os4G4Uz8BvRFeNCHuVB6
bJOX6+vGl+8W3yHuUa9ivNoGwlrV16/llnXmNj4zwlTwnbvv5MhjpQKTzWF7qUw9
Zts8LOAWNx0XmFIUFOF8TcIJih6ueyVbY3ATKtnVwfhkqly5bRnKbFBTVZZcIu0m
cR3WxxUvxOIWF3K9Cy683CHgVNqQqzTQZUBhs90wsuylM4WAAF51CNZhatF/Bey+
tAKMxNrbQ2L9zAeLILqW69EzzK+k+wB8T0CqHwdQoXG4lScpC8Pv6UbaQibuX8o5
iRBmXt+mdDN5SY9L5a3EDA+wdHQBlrV3loOtSCtnCHd8UllbEwDcs7n2RD+JQ+Wk
HY2ky6ApfroicyC+snfPGcV96BhQHoTHnwU5Xd0rvWyclcikuV8QRQhLxIzw27fz
I6kbGujy5M2B0Thvxjk4EUaFYRxnn6rfUUUxtAllc4FVyeoaNjrIRFu67+//qY4M
hyBSq1nlxH/jh6DWD8I68TZhE+3axq8V/FCrDAxsOEmX6xo9lFgrMLhX/TTIufpX
PkY0si/jjYZyOj5uYBanD2nknC3gnKVJ9ArsDF6OlmkLN6Od3XlkW5xk+vHM/9Qh
n5XL0/FaJxSwmGiAwe7fntyz/cJQvpvLvrgMmWhWOy/ZSKlyUCcUnJAOxb1LXTia
uzNjARdWD2dapYMgFgOeTfj0WWnVuvg6qhFC8eRpsbKW3nkvEYIKFBtcYib4SEMw
/HQIOHgFCFXjhErMIZNb1arbfcnUaLPdAVQVk08YKjLrMxEOQF6cKgsdbRJ/FBzV
UfgSNr0MV52G/qviwCy6pUH8I3incQBExTxDrBIa/f52B2evCEjh1jABu3EmR9S4
hejRiP0r8qnKYUKoshVYfRZwcGyOjfTN7nlk2m0SzPThSdDk2+w29eYhMsZkQEVF
xFM7t3LvizQ6n7/GEuAw4DW0u15S2lRvKdfj1ojmlYSMPRNiwuDF28yBpv1YRVt0
B4quhOOJ1GxbMSUwPLVmVkrlxk1e5zWh1m2/rZOKpYlr9V/C+WdwXhU+h1pbknXo
Kzsyt29FAnHdjWACjwkuSjSmoBhlri00cQfky4nz0PKbGrDoOgHAPrpsniajt4Jq
GiSbphDIghJFfkrTdYzG/aO9Y17jGd0GqJxxm5jh7m8w4/QjnlXV6gnG3HqBPgV2
osgTOuSLM/s4/Q4ojGTWV3iKFdT9rN9R5p1Xcy7LS/DB+dfWGiEd5Sc2LpXRQudr
11F7DMaR9pbqznq3yyLw/9yRwIg/SC0OypqmNi1sHzpRMdb8KNL8xTzy412ufjYC
HckZxkAVyFcw0oU9R42DHy6ZlNZwYMU8e4Rv37GCcnpfYqY3KBkt+MOGEKZU+J3t
X3LlpCpxKoQ9NPYZ2nwJUehDAdsRHClSW9tHTLQ6GsjDGyd9JrwZBABLv7weTc0E
Q5aReTgq08FepPK92O1VQAwpszz9mmuaOUfLbDM8JCH0yjTqk6HbQRAqMX9iDzrX
0csd010M71DZOzFwvAVE9ciOTeSrbaMf2tuIsp7U5GhAQu0yLqR6ZXxc4luIHpGd
B0hA8KWhf2LgwdVY8B0X2HWICO3Z2hBQ/RQQD7jSw7FQz79h69bafTumM7qPuWaQ
8Q1M1qJ9+oqnmWDAK0NyZrbvupwXPCQXb8nqmBa4rOVlUxEpfOZUwPZLaoAcl52E
1zhNJ0j0Jp+59E/5wu0RQpPJWS8es/3+y0flIHhMufDLV7H+ioupTI3qwjYYhyIh
ARehtibUG719/nZUrh85oRy9T30ZaCLchI70qAvBebGKgY7LFtZTk+nSMnb36n9u
/kiH4EArQYyfii7YW1/IewW2IpCDkC0g1YCZ8zSYiv0za5A5HntkyEI1tSTACwhf
1JhNAjNbHh67+t5C//5Z0tHYeRcQSgtP51xk+RbvqVNHTKAys5eiwxTPCbhgG+Qa
rQXjTlFuKTkuD9nwe330HY6QHQCR+XN1T9QpTcVbjRkawW9VGijNi896B/Zh6Nxs
iPZoebJEcjoDQ+ugKk5ajCskvCQ2E1C2kqWEYR3L9nusp7yblJ/G2s2nJSdufqtF
85Lafo/ldldQ/67X57q47Y8uzrWiRYDDZIpDoKkiAbhpqvVxzVYWWNDGxxPJ4pAp
lc0ROKTMpa8ChyTf/8xT9CIxix+csS8ZCpXSX1rvAwlmQ8QNCcdgs7/DEjd5syuv
0mZd/5jz/qadTjB8nIPkpPlOpjs5fpWlgSBD+u/3aa10y8JW0/dxPnldbI69UF0q
Do/Ptgk7QE7rJ0NXoauSyOurzYlZw4B/muZUx3b61XpPgg/4TNL1M7o5ytl63vaA
ZrVOxR98lMl2k+gfX6WG241OxSmKilGtAtze2nolDVGeh3pdUenXdhZxy+zXH9/2
wQUJP1DJBPuQSzerGHi6x2bYk2sWESioB9c4987Txr1lelzC8sZRFchV3TZBMV5P
Zk1UjwtAqrmu7L7EeQc5rIdXcfrpdoNJnViDaMsG2Nl9rDd2iKiSXDm5aQ+ESBWI
drNa/MZcz97TB+UohQA4KBECAuRAaIhZ3QQt7f9c7ZRhVLO0WSt1Nj2I4HX5Kl6n
qTJOwYiz4nuX5F4Df+p5BAzotWtNVBC75R5WuIf30JAguHjr542VKwv+Of5ZK/mK
mQK2nRNUK4XTMUzX5qjlG+MnDS4/+1V82HXKLjEkcVHZ4ybBw/Rt7/WbJShLPffl
HDLC5m3q0+nDr174P0csTDGf4Bg+q8SRmthW01396g2lKqp89ym9Vd+XhiiUr3Wd
hf7cWvnuSshROEDdh7rkE4XmoPQaaznPKq/eUC7PNbjP23wP1DqicotzCD9Lb424
hmIBlPVIdGkshlx7v4rGaWcmQZ8NBai6Oq4uwI3bVUnmIpQon6wEu8mM7najdedv
Yd866vCqMHJYoKbD94u2685tMoUdmHvgNxvuwFcCQaHIe3sW/0KhwLPUaTmKEY84
SmZx/dLTJM5/cn1fyVu9twe7IUP5RFacpR3+Nc+LboFZvT7swhAvT2kei/yVgl52
K8a9mHMuTiKaq9z6TpkRfKa8M8U/hYDpspOSAIINVK1+EVo34gKDBmk9MwiwuZJm
jYDZ2xN4HB7ib5x8nFmmFsPB1695cfyzqT6Rv7okC6mUSv8He47J7+3HbOGigmmb
+Z015UAccgta9mMgXXoWrqyEQ3YdTdneYeIop6TK/e4CG5oxqfA1uUA5LPpaZ9TS
ml52c/jWCY1kJD4RMq8d+cwkzwDGnl4uKvv4L2G0oZopvTla8q35sufsIaTD+d3m
kScWt0rMeyptbsHKBLtWmH+85107g8fSLmQ4caVj+Owzp0zp+uVcwn8FYZ6f+BuS
x1l2b2MWs1mOZ3E3NtofALk6I9oKoDFuGQLW4gPolRkd6ozkBZE9TtRPTEmC7J7c
Pl7+WDOJ75jJqDRoM3eQTurzRBR2v/RTPz0Z4dOgApxo6H5qR8NsCUdtvR8DNYCY
3mcnzvBjzNiuL6tQkxlDLI8qZioziBdMjnV7QISvCrIkzIAq/QSSSRDs4FlxYZrr
06kNet4JRJiR292W2vHunjMBC5Iy7kfJlqHPcrflUtqgX8XaHUt07pFwzGi2jNxj
APjKFIuM4H96BN+4BzuzqTKYuj4YzL3KwSvnrSxosJSrPf3vIT6CXmzcb8dQLHX0
by17ObOjaa8LuUTcJ9J63d1xAZMIDaMfNvH5NKrPLenrovXKNc0tsqW56e3wyBRf
5az8WtwxfHVBxsZ0IOlI7cEl0LWcBHzJbq3TANMmZgSfAGpad3mnG/iOzb3Wa4TT
Iozypn86iR8W8aAV4MusMpOfWwL97UmRB2aoiPNA/chEXnoFwvx8r44/+iJGfc03
HZpqfhKQF8aZNII84oIuUN4EwHS++RN7oKEHyJ4GKO0kEHzvyGNiL+mMku2u9v6r
+3Ok1igwsehxiGN1swPofBxyxBw+qAG+tx2jLjPvowdkEqWvlVmxEcgAG5kZHukd
YcZ4EDzQ4N3tRshY2k/WIYbbDoaW/pBkRbXPFyaYkURB6Jeqtj7E9Go/XLEuV+MF
7dLoaioQYXEnxmUNWO0p7F8rPez5OkJu2hsDpSd6h4PNsl2ZbmGiqT7DNYkpO87e
QfnEFt/+jR6oRUg9iOId7bBmDqAy51ukgiGoM2/Rs+UjCoycCkf5F7kgdeSGRVOk
P4l1bP7F33xyyEWZl/a4e/AAb2VB3dodFnj+IC1uEqNsnK7uWw/iyVYVDZjuSg+h
rbPlLHJuQOEaGpL8kyIZi5kM0PehUS3onM9jMdq9ZsrWTTjRojPUiQMrzkU6t+GB
eLAyg2mWZij4LAL/9U520k5IQSOCr8ykxUxNutXLykQUW3mD8UOkgvzAC1Bj8C52
AbnZBLEIISVbjJKphqX3ZWES99o0mJeEgm6Wao7I3Mu57JPpVzO10HT9kc4Jmo3k
8MnJ2Mz+Y3CrlOKoxxVwYlz8EDnR3yKjk6QaICzeBCiTK08nLzc6si5mN+JKq0P6
IoMDlYtsNcJg7h5QEsxk7J1WtBepjuJ/J4Dr3OhutcGm+e51peQdGQbhks9ntYg3
/efTdLcxXIx2ZLCScwUHJxN1AE3QgurTiG+VHB6q8IXEDdnqvTq8YeuUZrtt6TXz
VRzrM6x60BbXCXyb/wO+gFGvcH+fwiUSikzdsAb3xx7iV9dQaB5/jQRvPVtgZGaO
fxc1hlO0UgY4K0MEeN44t+sY3CXaz1v+TBELHNwvx+7Z+hrwUw7Nxl0rujbJkCz1
yikRhKCyXM9BGncTUUM9COrH01m+Q+LEi77bd7gADmM3T+dhzqA62Y9ConQ4Ze//
XAdcufx8dJqebMRAGETYcLYuQRl7CxKg8lYxNYCwX+jqYoP7E8j1Ijo8gI1Z+L08
PFSOvG2My6EC2BqDeOGEdpmMKQsqQcREcq62XSPo+LCP6zBWRIvQOIDH2QfP2IKl
EgWzoJXBYP1q6yEIYEcqD0EKq6G85YZhSD1b8gNzpYBCV6Vg6d0mOqueFxZdyNKn
fwjxhIs8cpoqPNl4SXkACim6znfkAvHUvOEG+1ZxcqY1YdEyVfmXSjHWlESTdwpB
unpRo5pwnKJhM0ks/XrZqKNapZSKDLE4G9wS3t9i4V+mszko7ZsZj4qVo8JbyQpQ
iXFQqu2Ca/Pa9rj5rnlgVm+ZKpbL9ovuNWhQnkpUgPt4dVSZpaAZz7pBKCsbWDB/
o65A/g7HUikA3RRT8B7YzSgfqIGmibNwaMZGr1fJaczeo7KQJAoNsAiCg+lYfLVc
tVBXEeoEZXeo+hcHGr0umDW7Mgi0AFybs7k+dBPKHWzBM0sJ0tKiqmHEZOTCVdE5
11oAxdNzamK5XpLLR8zVboSOn+ecLSO2GnUtnl82QtMMElqHaySRr8kj8a81sh9/
DV0ZS1s9LTufhSB6yb5TAcAvtRUzmg5xpVRCml4JuyOM5qo6cP856QB/4DYw0xTF
/z2XpGv+PA3PE0KcF+o2I8jrX7pMNp87sIjDxt2nAnE0IjgEfPYoueadUsh8cbf2
RFpR9k2HYJc55ycFZY0N+vp2Uif1il/KDoT8kpsKG3jTBFo33tCp1oo4afBtirRx
1yORCgGs8Mdz/VMtdJUcZrvAtzLq1ImJi30hsFsAkp8AfGBv+E5Zu0Hm3sbHkOQp
ERUSW/7fRY7cXBZy/RShYB866QpChKCPH0sdlR/g9p//Szmw5z5e53HU48IBmlFD
niRPWHwNiLunqQBS/Hcbm4b0e3RM9YSSGJIDfzqOUzjsdAkq57y/kIrm3w9+JBXU
W08DO3Z3cWjUcR0/9+bK3Qv/bmc30hSJy32Iu6FLHb/uhLeZBwBmefyQCBVHeEY6
tC72O6yaDBQRMQd6aouZdAHue6UM0w/sovz0iHPZsPoGJg3zKZKWiwUtn9nMvOcY
s11BK8lN8Dd4U2mcEUG8hd38iKCNZ3ksBlhywhrlBUu6L2N99eJr6RQhhKqgLEBe
1fUQ4CO9HetDXcz+1wv6KTnIb/b+s5ryzDCmwwmy36L1v3XcJrJv8Bhm4SKsnu5W
2/3xWQlx5C/hK/76DXDwlq2YnlE3cDBLtZ1aqTZ0mnW1FXHUdc9JsrTP2KNwvYgY
3LPPnc1mgLOljaBoHXiqE7qa9iMC981Ri1Y+rmSntsAxFrT96o00HTPLpzcaCxiJ
kbcqo199U4LzighQgH/6t3/1wqWNFbXJsCHo0F82ltv//R9/4dmrSXOPOxhDVvXY
VVj94ypp4VhIz2E9J1a0AJ3fIgcwSqVx+sQ9bmja4poO32fUpLsXdA1h09T4Jq8Q
yGISR77bND06mQhekMnYgke/WZFfFm4jd0tMdXtcvODfv+zytavH+XJt6FOT3tyg
EHn0x4dyVpo4sQOWFidzMFJD/DNdfQSUeCrZ+9KkIm5pOpgVYVmH8o+fXXfQNKYv
1R/VsWoX598vxd1YCsqlIZEn/Lvna1Tl5+sW6eGlb5aCt6Vl515bRjOwZcqr6ZZq
XIfMoVD0EVqRy9zuNaR/TQ3BmGLstqM+TswATpPDXVXkNnMgj8fHlGC91rrU1qNN
s/zjvd0HJVrhG/lkarsKZP45TYcPLgUWY20wNnRqogHDc13oP+elKfCHDaDbQ5pb
dp4zptjDYHcm/NbUp33AQfTSYHTUSwyICHEbbxcn4F6KkpAmuLpICpSJQiXrIfPP
jaEgr+AfItyTp0ihS8+F6POmMEZOfQxNSfewU1tprqTcEK8AH4fShzCQu1TeCdwc
OWKPrUtxypamJLC1e20Jw+oLrYWsP51aaj6L5X+bvvLvNZiGUED8SG5chmXNSJki
CYm/sW9WOg01RTwsfwEneYszB0wcp/cj+4iVuLEbOLekTFM29/MAwyjZsa1AHT21
BeXQ7PPjCUnpndBSsudjJRH4RKyGhz2+hj8+7J1HUOd9sm/Ii29dLL1nSomOxFm+
dCvGmFYX9um7Y4BYr/DXXpuem91FjVgok8HcuSDONuFDzWHniBBoBCeFG7jfoCLb
r5yAr2EqF/Z49b7mCPhE2pH84jMHN+CfoD5tea7qJBH2rQX3oefyIG2rf9PWdTZZ
ISO8kY/y2nyezQzLrEqGFpoOs/anzif1SNQEXTYc2u37RoJnKibAeBje5oVJwNal
DexZknDW8YJqdyUkg9squ2dz4031Nyjm66jjdsb/7vaLVCjNN1IJWchNZPB1u0tZ
f3nLriKrqXe0MSIDqvtuVsS5ar799dLS+Wa2kQZm0O+adT1+JTx5XohF68W01k8K
Y1cevob8nN+XVGPrw4eBncfYsTC3Jkk6zjb0apNBhzRmV5uIvom8P9FzH6n63ONU
6QlPmmBqK/aqKIPpXtjsKtWiFcDwY9XRM59ymzXpMXcTS2oWdvyPKpDBgxT2wV1M
SLtQ2VGuGPSp8LV9dQe+yuD7Ho5t5Bu3tzO3u2bMKhOYbQ7wfK8GHMmSTLjKuN+8
wNbjiZcaodXaM7DPJSF+Qx2oFg38WISLztWXWeLccGTE6dPwvZSSdGPvMIyTlV+E
bX4b/PzQ32pyNuTKl7Xn1Zca/mmiuwE1H62BK78vfX0hGeJgVdhzNXr7n1SkUQ23
8N7U2Ge+b5egYEfu7RD02Bi8tvyBiDRFL7x1Cl83ObOX7y1LHSxEB2bGTPqfaBBw
nrrxytOQe9xfWxaTE0VEyP0bMIiJ1LK5yBikeD92N26nutWI1ihq2aij/L3JhL6o
lXwUOuUnwJkpgOgA/NWtpvQuVHEALy1CkKw1uGidStx56tB7MBPxxS/KlAsfmlSp
fjdQktZ3QJ20gvSds1eGCMJqDwwEDPGrMBtH6YSgRBo6XWc84WY1/dU0a1psQ+Ts
lBh7l+K75VjVjsJ4mVfHMl1ihHweKwd5veNodfE4Zmq5qLxqwDsVdA7Z+cKvosOi
KtthLXrAtn62p0RAtrnTFTJrf+2CXaE9wiWNoGjd1FMzzxMq2BGM+ep+SzQHkW/5
bBOY0EPiNaWYzS9AqvqoAjoJ3HgvvBH630ERjQU5y/LjnVTfj+Fm0ylQU7VMhSkD
2OFZbp1FuQmP79jYJoaA+vFR9C0ZejgOKGB6fHzMxOa+iWNzcXqQgqnIQ6S+4qEI
yGQIzMMLz5M6FaQk0YOW2dvy7FoORjYdPELN9ItaMRO/ZaeoRZi34sVTUT5UYmr/
G9dLnNiJyn+TL3RoD6eICh50gSBqgX8PKYvqho5txsCM10xaJPX0R4Aj5SkB2Nxd
b+3jloCluHc9SP1bxcLYYZ6T8uPKWuI7HBiOI2qSb5WLf8g6BSENdaX6XS9dwma/
ttON8u/X+2WsgcdVgSqaj+1vYFZuyJ1LB9hSzLz2whwSYmAkBbOhfLBwZCnQoXER
BzEZKTihW48b/6Nl6pYDtkSTxQk/M3YMV1DSEqMxLowGhH+iA5GwDN3Z/S1ipOX1
aGecpcSTWgOR23AkN+gT/Frk4QTaO1RYuIxyM4E074w6SAiNs1g8wmLArF0/ircH
UpaPorAAMFUgh3NZzKY7yZJhE1duuSWort7sFUW+x1GrmyN9mihP2MxeYISNBUgp
exJgJWJuPkEfqpxh1Y37KmYeKVmMsErXwYJpuCPo4wQHXD+TZbhTzAfUVvJajTco
Ao5vCvvMbgtGoyXZwTQCikfD+3/s2EUl6SIb3vOncVLu1x0M0u+8Ni+4G9GVlEEa
BzMPfhyppiC6PgW0Wef5meP9O3EVgVj83YIDn3doKRwUUzccJyC+wWQMkriEnxgi
6G6AaYp0ymTjn3PeLKeG4lrorWe1bPyiix4TNxw7MrwiCiB8bryhbNnggQ5IA+Nh
lI5VjRHxd56aef41ae7cPmOOeHteSYyR0EoY6wsdmJnfXmWAPq2YKrZnkqPOz077
1zUAeBpNiSnHnoNcGgZP2uY3neeWZP2C4gb2+Ee+WsepxxYvhWN05UOcZO9GlHBu
oY18xT8YYj4rCA9+m2mE49Ym3RDCtGzw3MOt5aigkQV9jTrwj98BcAQMYITwHBed
s2AqMpnSobz6TGMTHARIBOy1tScGeic4QgWH80hNKJH6UtvshAdY1EtpRApy0hs3
VzALIaCg+QGFDtvRQVXX8jMuWT3t3rDEGwxVvlkX24PJvglCGP/ALfIEDWGLxskK
4eEQk8Wdx03TE9G9hI3FzSmGtkCK9phjVnYLhKIIPsqp63P1bIlXaOkExyx7BIj9
3UitVO+SOYa8O4pgjS4WaqmBgpRvSrfR7EW2GJ6DV8Y3PivGWrUACNtY79KunPOO
j9D/6YBE7ndGr/VgNAndrfPNzJbSQYvEAmcIH+WCx3y8ptGdFNXmrivRrZXOdgqx
x81+AxdJWEHQUxfigI9zi1fabsdKTEG5kJteedFCDiA2mFeYelzWtBwNcbsGipQo
BkYxWFsoqMst4ydbJqy6RO9dxmgOVlUa+C6fbMp1uWI8CvBqTLFJ07OwzaVHJaSp
Fmm7oGQn2dwYeiaypr7r7FtC3YpDPky7ed3W0oH2XoELOOUfVkSK2nVlIlRyoKht
MPaTXL9Fw1/YzLOYYGgl2mGnrQtL5x05v5gAvPMQcCxno21t1iJpsjwsDPRzqNMk
nRD57Yw65PfuKiL4LxRmNYGEIOzpMcOt5tIAB7BSEPVoG+KzdsLvyT6o9NZMZ4dH
K9dcEVlrn0YcUZt9n3Me9m5k6WJWqL08ZwASyCj9Xvn9tpuK0y53rju2YfQCHCem
EsJJiY0cJl55aQcnaKl0LbbWf84HNC6bpBv2mt/9tsyGg1CshA2lPGJQdB84+3Ia
x+1wxzITt45G6tdYboeaOoU5qqlsyinsRwZRypWO/Mw65Xn6D3IR54VbqEyEHQ4L
M+t4GYoiGbWV8ArC+p4COr7wgNJk/uglzSBKIlwmCmOIrxT/BfUpJ7bt/R2wei2e
MIzKlPUFtBtbUEAHuUCr+Lk2+q8A0biLvpehVdVCM0eo2eX9cQWnwV76HIrPxsXP
T2fPxzk1Ny5cexPRCVyah3dMSbdfTS59YtiJqGMhCryIx9QcDVYyxkWGOMy/hYEz
14MKlsptzNyXeHhEeqCAWi84JBZA6t2VybfVl1Q8StlkuRSx75g5utCPrkycX5os
SnPOFHapeXPF5HaWpOVIarVRVrUrHbLcVrk+IvHSRztrQHg1JUGnkGlB6XTC10mQ
Oxy/xxnTc/Nn8PgqRIS5hY6PfSYdLmX+v6iGdjaajx/mqSlK8QDPyeDV2p/GbqIH
MaIoxL5C6MtgJ1BXL4B9cKH3sInrm1qpkJhl4whmLt73cQF80r9kwcUVBe2IVD/+
NCvPxcBgEpsjADzcv4krB5bH6BM1eXyMSXrUKRUvRYsiN/ZDo2wGEPuVIzDZMV2g
xOy+4w5H/IJS4LwJE3/FaK2Hb39hFqo7/XwRbRFw2R33tn4JRgmEgpr68CRDwR82
lGUkHioSC9D3B7YgI4DzjoloXDfNY9fRw13n1NW9bda0AK9GuVaBkHR9j6pvNxxL
TUt0adBb1tDJq/dhrrm68lcXXBQ6DbmE7qlKlk9hoTdNBh4xa80+UFLgICdrCmx+
KNXI3YMsNSjGQ+3rLUhKUHaESJfmWM5O4tehh6DYW8nA/xXdE7gXL1Pqz9xw4neD
JtBiH1Lz9NAimopIt73RHh80UA0uKASPaAXowXZGQPmH84gAHDlYN2iKz3GwywLe
bKqB7dEqYY/h3mhkVxOwrkn9+dfx1KcI9wXXY2K9ElG/NqSdgj2kL4SpltBSlU3q
pnXw1fB29HrFvMPBNTaUtchQRLdMl0QoNr40R0IOTasPl1eFq/SrnQiT2z87C05/
HybL0fTwtw1SJfoNM3tXvDIXobifVbVWMFgtWhb1RamnQdwVx2vBpx9eNfcQ902X
TZ9wZKkKO2galDKFbwJBldktFrQwWAKxnpZjIhD3zhhbbSp6Kx7PN+y8DtXsdbq/
BvjdUcom2oyyERYomjj097xq4mLMhXpOvBv8xfwYCn2saz24+qhZkpzKJEKDw1bk
BjalXYkyVfkeN2WEsNLF1XiD+ESMNj+dIlgvFvO7XZm0lBUelhpOY2qWCxSP6TIU
O1rHgv9dq+jm0CWd3fAdoIYz61JtIqZrzaINbhPVqE7QSDr1H2QgZFtYeVXvw4p8
p2IVp7G5i9D0qCRfH3Zi4LoQAM8sN61rNRAsCSeYv5dAOez4Iotu36L0VKwU546o
FbLbO172AIT5+xerrqYA5Y2Z0SCdIpUsCPYKcHrRE4vElxcwzhR6F++/9XDje0iY
qwylWDo6QSwhONc5tKo0BE0HDEPJxvQz4T82gh0PfXbAcw3nkHOvKiBzVBURpQF2
bf3jTr077PKESOwo5jBiowqsK9KVbWdICgE3lLPQ6Y1SDWdJ5+Kz3hcfuqgzWDhS
agifCi7vgZgtmTP4XEzEmgy72PGBryOqHTLN4erENA3f86wH1mJidrdLHdS1UJNf
HtnJ/C2E4JOEWtw2SKyRBqoeDIW7HodM+X35nt9efzmLITEfBNgXN8dWyprvLBYi
z2iXUWz67m7LE2e9WhtWfMXGrX0fOPHsLUaAoDd15pGvPsikewxu1VZZPCM4MfhZ
2sMjHd2Yt+lT063q2XEtN9CVHV7QPYf47tyHWOvBptpNj6kosDgHGLPZtSt94Uao
HWgws+H57Xc0bC/wCuX3PvYSMCYU9IHe6SPEMPKGuyCK0DwR89JURprYSY7Z0TWU
cLoZLXNhAmBUR3ieawfEo1QmhUI9w+0wGL7rS2zeKIy/8x/T+sUg7De15ebA4mBz
5cLPPRdgGF8lmmnoDKGbA0MQtBNXwE1LRRmJ1VtK/pKh2aeNvpjW7+NsU3P4RpEi
1ZiVW7Ch7N+vnQnABBR92UwrS+vMfGs47Cw60aOSZwaMH8FVM3CJfV4ptj5wfm33
KyI43vsKKhxPAycr4whdHwYyix8DNMl8ntTZnip8DpDhMrgCh4bEff134yq9h5jj
DfqOMJe77VqhQAOxTN5NRFN72zqp3ndHsw8dZqHxc7mvRrVrQtuTPeI8jtlER8t3
2h1yzItkQBkifhYkGnh4emd4esStSLjjGlETxtJVBJMzI+QiQMytGlTxdfgyPpM8
7vPlbpF3vZeP7nJeGO4dFmaw1WQ2gx3E7ZBCyxIVuQbHYpE73GduWgjHeowr3r8z
/H5WedZ9EOlVfi4AjXNaKnmdU5tr3iKGoviR1AoqiB4j312oAT0Bcv71GqUpMoQF
g/bpyrMc27ooeX9W3WYlodLeEGYPC0jFokLF/aHW6bCsNWL0YSTvdfzRtYKtplp3
AvZGY9A0I4e4f/xPetLg472kNQwbEVLOVIVVACeFUqy9bDFgrqy5oINXtjGiBSPn
8M+jaiRGeo4ntYn7YDcPGlkI6kjk+h10mZfUmQ+8btqRNwzU/AyZ88CWfu7kaDee
e+gZ3UILWHCYrwSP4kNWStP7oBRO8wHslyDNAvx2I/tOLeaZG7WSgiOvri5UgAKM
uPUO/1P6PNOotYXMsik9V+B+c3BIwiMZnXitqRpBVAVNYYpXR1gYwgr5iAVsrGYq
KqPCAR5ZFkgnKE70Ka7luNKK7y7QA6RsNoxCP/jXvGjID8eZFhKAvKfotSQjsUbQ
/Ra5w4KAiPTzulCxKLymjIwLDW+uVJOSiy0dvTbAvunmBv6lX/GyzjwDErRkjqLl
/Zlx1FKZrqS56l7bEp0MdfatvZAgRy6VNWqy6ClD9te7EBjMJe4qaMj2c7KZJVS3
2++K0P4G9TciknjzxVuuMOfxbWe+l6FNBwX6Qb44Q1vYNmm6b+Dd78Qzp2Rw0mgW
q07H9kzLlGt0dpRkcEcubKLYAjvNntTCkJB6XC6nFJYU67+aPDsffxBBFp3FP7l8
ZXV6FTdL8OJPkVk+7N54p0ol0MX2dnSAL7bEkJe7NCq4q7jLwJiskWi2PvtJpSlP
2LHD81zoLkjG+D17TPFLPokUlf8CsDfCUhkeMugknQXfRRbaeOtEh0zH4wTz8u3Y
QpirCGc809P3UBJonKK7dRYM4np0k+BmdszmhewWm7GLFvMopF/ksW+cJQuLoR3E
BzOgbqPPkTdTuMciJPu19yVyPGTW6mYtOdqiObcsG58ZmlZk1BTVonmTI/zveUoC
bypqxGx1b7Mfq2s6wmbFHsKGHmXH2PIgP+OR5rbfJQJIQAXda0ENaUi1dQD+yCnW
PsqFJSj4d4CNEzbfHDM/o9IiFX1xZYstviys5GNNvbbt9hGpTXa+Z4VGodM3CIP2
6vxE/j69r/ki40Ks/35nZDmd7P4L5CC7b+8RU1f+f8qIsgdajcB81KT6L0QIMR7O
TNTvjVYwzDchbnlubB2wPAYnZrKzITLWUtwkgdQKzHyw2Lvv+KGkg15HKmNuNMrd
wQEGJqpU9kgCTZnDforGangXjU4ilkNhs1Izyhv8wAoSjd74rdh36CDmMJzuzMg4
0U7hzLVekpsdMvb+mfzkglU35loHUj2IhA1/Ydapc/PWc2FWIa8bxxpHIrK/YhkG
pxIEFJtdoCWcPMLrB1HPAfByf8DQYZ0PnsWxX02eULRCTDvqVM65qzNDfM9PU+uE
zH281trK+0a17fK7LtXTu7C0FAqozzfqfQnIfuOU0MQ7VZuulV5RmREhXfx/EmsN
fMWStPpzhiY9BjlLlomQ75KkV8XNTb925115hLDlCqHX70PLC/fvK3B2mIz2Hlm/
0b6WkvFnllKN8gtrXgzj/txAMQ1CT8yyi1Ot8k39wtyPj0C148HfBr4SOQ7guDGk
4DNQ5nh4vqyx+iCry6szfAXf6+U0uzbhtbcKT+vkGEDRM8FTabQSp4ceq2QcYLxU
v1NVOk3ZehvbkvsfK/QNO8nwB1QfHzsLBXgA9Fq1uQBgGjuOZcFH1N+WRst/TWQc
RxaZHvTA7V2cs0Fl6QosMcdJVV4qG9SP7i7vryjQd44iN8GTdwWUc+oS61abzB1D
eFCT9Ip/c3OFtJqiZJSvC4X5TVvyhu+Pn2C/dmFDJ97kSjXvTvXR/dUiVbutwq5B
7Hv3JVckNRaclG8QearjJHVsD0KWPQfKJ/HDZUDcS1CMNx7mXNIwGHzr1fRTrfpv
3Uj/+xHgU3lZTDNMJLlT0P9s/LZRYvaQyN3hxnocbpPBwTPc/SjwhMlvFgHo7tea
lF/aJ2UfAAzUyuML+7UxIobAjbFGPAZhUjLZ39dpyzKFqU4TspbhMlwnqgVip8Ex
dnTAxugJfCqZakAUBf9OGiV0zUfCuSEERWsd9Xp1b+9EyNwC8m9/NlDNIvmKjqYz
c0udGfdsQRZrF6IRdFdyVKKavGIYTM3KNfYlbanIIXKNBgwE14CKm9QZFpSluD8p
xbKB4n2TwIgGG9d0PsDfnYk9ALeCqoM3tBy7XwhSi5p64GePKIXRrudFLFqM/gui
W6tTmMvFGu9w5oFI7/RBTAeyWZLgjcjcXqjGo7WmoluOotstXBG+OcAW9N2JEanl
eiHnGj24BNM8WqSsqNaccV5YICsev3TLr1S/jOSjQp71a2jcsjqzfmW201EbqPqt
Y5yuQJHgetP4qPmGSzgC48OrPUsetj8Ogwuk2X9djfYbbVdtuwYpQHUp11afC/Ba
y3jjowxe+GqTVX9GbjVHyRZKdeER1S979vsbpyw/mHXnNLDD2oLWmKzqhpKqaI/4
zZUB7huwYVOTngttk7dpBt2qukShx8gakLxi3WKve8E8LI436hN8HtBWVRUJpHgT
3Ar3Vz3NXRjQoX6ja+SEQkmVbK7WQEv6XpE9Y7iZVo3D8PevyLzHlgxGtI4w5kmd
IpVIv6od4lLr1HTZrn64LR0kIDOzv9ux5fGxSwABk5mYnhAkD8AG5CDkYPVnlZRy
Fr064tRDh6a7YrwCQ0sOdjhyEfkgHn1y07FDKKjpNxwW+vzn2B+7HSM+fMnFNXWy
ArpEIDHYh6sPu8fH4lzD2QRI1LIyi6d6+jC/yZE8GQpsVEv4fXCnxWo8Baisiyf/
DJUzJ7YUCRI4muFGWepFaWBInGFpADsntX9tQBnSKRmcuKsYC6YaRCeqW92rl+7J
8oATIKRnbXnrHqbu1AO7W5ZboVwflaa+exIZgNip/4KMKsNToC7pUIXBR1bqW6Lz
QaLDOm1+ftXmD7dNET+DYMtQWUeHl7vKQ28IBxqxbYh589cROP+dvzzodJ5n1Alu
YxefqMwaqKKMvzJEN67PJ0UXIzfNDrzQpUlFlmilyha+SdcxTXlczL1b6o11Rkfp
PejcPf84jlCyfmvAqqIG39mxYLDBXVHn1ibYOQhNuWoZi2tXrgwQEYyLzUFahXAW
ERszAZ1gzTfjayVNMGJ7oghEdkAYtYZmRV3aAAoH2sS1ANJtcpsI4WPMD+/uRA0H
iEDBUZFZzXqJRW62i/GPSxQuFISRMQ4tyNfSsUk60bXrPWBF2ilHXGSDagAhU+d0
OB6+S/kaQ0ALjgeN43hu2J46/lehX9XCht5E9GEqLbqvn2237jlQRdTooyQFceFR
N4QPkuPFD3v6R3oL6PSlxjfZR1BtT/XUN9lb5AlMEtPOYJ1GhHYTYLoImc8F6ya6
JuND0P1nJUbwp/a9fd4GN3zcXkLI1+mZefL0d455SfcJoxlkYFiBaCLk7FQfHXBT
3TejnzKz4bouq78g45+EG6A3gn3ck3zJFpnhI1Iceyc/IAkrg8LnFZNkrm+2Zi1H
HpEip5OEbEgI5ey2g4SORSrlnVkeU33SWncgNtNiyeutIwSHch7hPe/SQwJPm+QK
TtHsop39au52gznoyO6oreb+5/r9cV2ZF2N+1LNClwEUE4mDJsaG6SuKT+J9P4PI
LyQbCqQjEvggbnJhVmH4RvSnoCmvebCr2oBwKiiEgdwCEdc6CxZ/X9n6hV5SBRYA
D8XWLKZOpUjO9y72S6LrwDy6bJNbrOdAye+EEFDeO7yZ6o6i35kJFDsrs6NkCesp
tZz5Rika42Halz8wBIqTiYg2P4SWQW1hKXC5RwfaU5ApDcwb49Xujmfxy9ava177
s6LSmCzzhB0wdMVxSiim3SlMjw/T6FJMxodbQEnh+lVqEe/vLlhbdyFvb3rIzNQ6
g7byKvr4yYFDuzoYInzxe9LBvduNkyrZnL1d34BEehmtQ7v7+yOf5mBXPeVFiRVX
0cf4a9qTqNswqKL4SYpXyrSJBDqdqkeCiGlmVF/1Eq8yKuV12vk7W/1OVHyTZzum
8MCUM3rn6Kg+krUVkiC71X6zQrZWPha1lF2uJzJd/aU7/pVHQBNTs/7wZNL16CQY
ZKIpqNdTySOyLhAM6uZb+9YO51f7MsWBC+QIkQsBx00IIlRatlWpYHFpwTMxjn2T
atVGJXnmkO0FzOLnI14QZ1GLjBXQDfDi9hxE6DjGTgLJbCvssimLUsuT2rW9+QyO
GL9K3JRmGbBPQuLHVV5WAYEtGxLYlmSSN5r219y3hDFcX07D+itQuXpEO54qZIIA
+zA2tOnE04vNw88zFAcX9b9S1FmtM6Twcja9dzXbMXUZggqWcNNlHcChGzay+GDg
TL5j5f9uTEH9GKmgWqjre1ZiciPFomNFeCAAx5DEQpl79RCKKMg3s8txdqZo9KMc
y19ZmbaO9saAGivrW8rmJL2M4yAiC7m2QTUBKMPcD8dz0kIjiBHJKMrMLt/GY5m7
JxQA73dYQ+zsN20GU/lmQS/udh6Q7ysMRaSWTe2pD4K8nlh+JXXT3wjWQh2upz1U
YQ56ORB89Tjq9U7sNrngnPg3f/eEvXNdJZJkSodgIC6uJ53MSv+1vEt1tGDcbShP
F8RPW2EGl1Zzgte7Yxex7Jm8AhILWkbRgt2qo8XD5TzAP/i8vVBlpvooBEPyYRnN
Q6KYDOvoZsVoHjA7kBIxAedVLuj1oltHETUzMqmMvLfTg53cQJYEF5Cqjrv9CPAs
r9lUnc3p/4I1v9J3WN/Nze/NCFtt64GcvKUKSlGWDwmQlCU7WKxHqDgnnn4sW8yG
iR0esMsrC0hCqUhNLULyRAZeD12pLzbq32PKU3otXjotUT3tVSDrlJ8lJTlgnWOk
c2jg2ZR1yoQ2hMT0smdeyvVUtaTzBnJZlX0BVEYqGAs09ViVb/S0WryHKAMq6Law
nTE3Jjqvs7IaCPGq7bVrdAXifhp86GXnDdAZhhN/Z0UcMvE+khQvNst4XQ16Wag8
pXuWbEY/5C2KCtqi7DobG/2q3kO//AbEXrgzg3N11a7XM+y4/icVbkDwh0FC4MW9
3+XRcnRqebyQD78ZXVD7vODi4xIxPnTuo/iAp6EeIKQZA4V2tI+GB2UiCuc2W01W
DzaBbbdkO3PhO77QeLdLpuBIyD0Qy9L9gqLOQAwCBXAjsxiM812lfpPRueUuNAkV
XyHakGJbhXKZ6uWC3zdYgIWTGYe/QuWiVAbnsmAqUG1uCb3k4xyuMOBYUPLU38mZ
rkSgi2P18mQBT2QraJxo+TvwPw64B4n7HXvKuIr/cK9HHFHg+zZq9Kmbrr7YPfj+
it8sUHyOofOcNzcqOZKeKdUHp9REtA0EKMIqINuJ3exlC7hFsoZNfKgYnXwExjIS
/fAIXWJAdTmMQSzBu8fQb7JtIVWFhQnHoFSxRtdphTXwNv+/npkOkeyiH6ntVlgK
BL8CPIlFwyhrvr9yfRpcLOjnYJbiWiWJnRMu9dSIXkvMeWa61AaLYAp1wmjo4gmy
LI1CuzWJmaguw6V+XNjgSGix3AE8s6J4KQJ91XZQQXLhqxvyECOY1HOer9OKfucE
q+djBm33HXtFv5JNmZtQOpe0UfXWfoXYNnQccemnXiva91PuzCT8sar7pXzY7UW3
cUb8D0bZ8ZtiTzzQmZmdKbz5bg8Bye9qi4ceiG3xld1o7jJZ4e4lNhD+AEv4YTQF
B7o7uRomZdJFYz+eSypbzwZD/X5OOWui38aRAq4Mpj3iLYOYvGwqc1tWVp3VjH0v
eJcFckwrLM4J480WuFx1pESEfVpJQ7iRq3mwPdymHfmYXnqd4SwUULEqV6aUUDHL
1YENU17byMwPMdCshqMRaBq1uEyCb+slkpW6zfF2Bmq/FvJEQ2i2bQ+p1Hntp+ei
9nSoczshHSALL7hZFosPhfbIu6u0MOIJAlg1xtMOLkjVUQtm3NeQrGx70eCg1B+Z
ku6NEWwkCijNZCazh2KA9qDDLlEjKLBzA3YuUsm5wJ1awO4p64lGoSdRNx5sMS74
nhC8kQBKcXdQ2Hrb3gky15cGi+qOaJ6TB4bPVeCAzqw07mcuurr4PTqEyZSiWrDF
psg+g9DRTj+gUfRq3zdXNftcqWrdspjpJ17tA0c7iKn7HnY/BWmjKJbo4YoLZ9I5
HOwbmebJCJw4JaXXfPEUMcd2EcgmmAtwQxEgqz2TdQL+mnOyWGf7qDK4jQDkGAPu
Dvieo77UZ/RvkpNONAhsuXPeO9rzT29oPVMCr37tQuGspPPJQKtvSOfkXIZx34Zg
QqpQU+VbA/VfcayAYnucWBt/qn9Hx+/hsL8c1D4ZZOOWX4npm/kMEfr7ivxEtWxD
qjgJbRax6uNQL8uZ1rrC5SgrtbjKS1rdzHRK0z2nURa7G+fjVpc6AcY51EYHOOXd
EIdv3petbzab+kmWHWzH6Okeou+CIgDp/gpKQ+pJyS40S2PzAJma9xFphORB3zwr
PblWfApmbv37VhiX/HqUPLj14dFMV8f2M7B2Ce/nwXO6HqJV7Hh79CTNcWCB7NUG
LzDkJSmhjrnr2ZwYDB+pLb+BwG42XQ7CJ5aJ6hUGMUO0JnYdwXaPE/+vrmVV23pH
/7OEtH0o+yZIWuIgyQHMyziVKCkUclQNU6qQBc35WIV13MrAmgSd8/ZFAVuRyU7P
fLjkD07YO4m6gkj1mRqmoiX9cxhyrVvEMkOC7cOr+gCZ2Z0T74kNJjFdfVIDWxjl
77KWHzEifrqhyonSZj2uva9eJ5uiJxw2KsJLEEdrd/yRth/GGAFD6jMsLLPXFtOg
ypoqesr1ogqnfu6fpOoJHTr1cBwTRjSzKGFrD5nutm4b6MdD+fNFsUDSGJdNadzY
9hwHeqUswEDCEgP2lZ3ddzLmSEb1mRVgAXT0sHuTbsGvkkW8Y50WIH/dZ0FcVtRQ
HLqfreyjwXutSRxNKFq6EenfDIAWu2dC52T6ap8xAvSVBW2o94gJXbCtg9dtLidk
DKWU5LgpQmTNTV4m1aOWau24tyc6AZI+pcxSmii8GC8F9gBlaGIHzetUX0PKqy48
5XBC6oiTuQRO+YcGOkpNv9Rfbfjyz0FfEzaNAY0ulRZBc1KZk9vvwjtGv/lWo25V
6dbxu2TFGOe2/iz44zqSYwhtr6RywemCeJ/2NO0wzbOqbFCGk9ZTSMNMeWa4/4cM
v0OpQCoSnY6Mml6yumf7UdTBHGzH/9afjtzhwTf5nga7QAXPFhCToKn4X8xxX2/x
gCL3SNPZQoH65YIP9bHQ5lfngfDBnHzUHblC2rxY2V8D0tVkqtsPOxxdlbkmI1TQ
lXfR0b5d0MEvk3Lrh26QwUNoQlAqvBaj3fgletnoeB8/P/dbLLUmIq2QAVldYiLq
/MygM2laz8oiMhtpJCytt0wRYI8OP/NiehVrCWsJihUpijDz8znhK6aWvK6KfW1o
D8QO7YVaV29k6gSEQ5rMh0mnkyCuvhTs9CMrKeKk9V76HL0xxwkzv2dlAEtmfPOf
0PDf/LlcJpLbUo8CmDX/ivbL/iYMwcZjSQq9/13EIhWBwLwoGKatgr5avxrJnJgs
2amnDyLvneeNaQ6JjmRUvmKOsbdDQ7/n0WSxm6Nr7eCGIe8CvQppMrmcwoPT8Aoy
q/CY9kFGS1IjsKVRgf756xVra/hKeopeEqywY3s5U1WDuW8qrd7QXtr/XshWOuyJ
5NM1sAKyAWXQDzoml5aUatRxHDb6B8jE1sLf7sBEFJdcnxM9EfreYypwHwGasb0N
y+BBKgIV0sbO1IshAto56PvTVnm78vv5EmUjacYAOQpVfUztRlENEYDRR/C71Fah
w+BRqDRFsH0C+xeh9Yp6zEUSA3Sztf9Zj2yeOk3gidB/8lcAfNbjsXgoN0XDsnV6
pSklsWeYygkbcEoywk3biIzZ3bvQ+JPJgFs5hxWkeJFbKqRjF6V8W37v9jj5trZr
Xgr4oZPK3Je7L+fu/SjJ4Xit0c+RtXugqFFCUn+ND3qXhJySw8HDsB9/NXI2s15G
55hiho5/ewFYB9Dg3jmi5/FlEXh7MAuCq0m4ahM80E3S4qY20o4foUvaEkTDsD36
kgSrjpSWwWnc8rMQuyFiJBTC/luTtnkOlist86NX9b+etHsaMHJnBD/SjvMpZgUy
VzxJkEB6+5M5VA4+oGZhH2H5Mpxpb8LkaElxY/MO9tkziEafqpdRjXhEJ9s3Sfam
MdmIwokFu+TfNrWf4PT5GBzYMwdsNgH5ZDu8nw4TVO5/7raVRDoGrSk2XF2EW3Tk
LSWlVL0bq4zg5OwYkUHljwKa1uu1OU8HKSczcka3MqsCBbilKhNMGBqnPfwjGYfH
iNHaYH+HaUbisdt/38T+Mw65ACgWvYMND598GupY59I0uw3klgHU7QE6z0uVBU+M
tHXOF/3pnZqxZobDVAeL4AuO4NUGdDGZp1PYEHKPmcvh2uaLiJzq0PwUJl7SXDB6
gkki5SSIrTifdgVzjogE6pkQExySRitzqQlIfjKQpj9LErMRjMR8RLeBaPdqCCL4
32rWaEwQddTGf3MKATPEaFe5DQxdwgJ+bqomftWXMtZtosZH5lgxETQOy57p6GaA
EcC/hkYwsUPuzPp/BCCnN2Y6A2lm+KzZuE7hxm5Y7rYH/NTUO+na6U5b51zhlktf
E1iZPTfaxkcDm12PP8wO6vtnt87BtxjQsXotRDiWjb5LTYBEjJLkCq27UyE8O9cb
dGvBobU+TI3gFy36vtpUbNR9rX2M/7s+UyiBtj2JadYCrOyBxvCQs4r4yFRAcxXh
M7L/dLixHBr+oSE1QqLzbMTz1yIN8BgA+jdh6R/A1+ZW9FmgX48HLXUh+EayT/Zk
kxdf2sk5mGKPvm3bi8WwNI1+VuULCUmtSfVFS/hOSWC4SUknvfX+jFQUR2uh2N4y
Bf/X5WCfsedNuHjbFpmI2swVtVgWQHfNU/yik7dwNDJJ9QHq7XfKzCoowLSHwidY
ooXHWZ2u4av0tbwJlH4aIqd94Yj3lQEJSET9WXLv9FH59MPlMplmqbRfqp/qdltt
soE7eR+/XyMuykbSw7joLPe3379M8ohoqUPpiTUy5kX3b6xCuQwzREy9aOmE8B7t
UBR52apYCWQO24dgUPVoVeRuNixYYaib3Y/L/5TEePQPn8q60TPNG4T8O9weShY4
HD6csFpotrGAImpzBWthrPiWgSyhjd9/ueY8j3J2wZdx8tUyIwkIYEPASq6rnnSv
mV1Ax5Zp8rAvJoDQ1h9OF9+xY4TlkHX09ira0dWwp/3SZWGS5G+638j3W920rAkl
RZWpZOCVFvmnjqFWHl2rHizaQ1FoUEbKF4mwk37nE/T6jkfy2Wnc2oi6/U46aT3K
musELM3MzL312Cn2XIqIMQSvYBqWoPJRG4hgxU84SmTn5UYOObLVf7YTU54pyqxh
3TFCyzKt720tTHN23us3VKPOxtqm2r/D7TiCgYCL+BPTmz5vGrBNOp3qPALylQe4
PQ7A/tmc92+aKJ45lwdkEXgaTp5EzasSDWKbe8XWdG2uDAAQe4eOfIbHPs2RWj0s
igvrCJZniudSRr5zVR/uGoT0fQEmwC2ir8xEaAjKxZVanzt7yqDkxPQ4SXbJSrGy
ATDgzxRyVPyw6touTDajn7laXLlfmf+a6cswIItAQDc6iHfdfsScwh6smAysUm47
DK5zhwiVVMVxjZ05szoSAkl9EAPXN9RbsMII59xfgBEgnIRoWfyOgIFqN9oseUwd
hVD6gOAHZcqAEQvh8wkfR55xEjzTQKEYhDPtlaM6aBg2lfqrrDPWHLbspxmIhOFK
+MAUdC4c98X1uOIF+0vxUc/iwUjudLoDtBLc1X/DljGoZOxi0CzGGfU5UH9OtYN+
IBtEJzYZuOD8/dpbXrVJy8D3gJ9++14M9T4YvZg/dFyVBZxnO1on2f4Ib9WVUisK
73Ya7Sw7w+qGyokfFDsj5X6WnY3JGr4suxTh7NfiYjo4KU4hAxSGw1RQ99DYJnvf
iGm7attEdD3e3CKlSLp/34tDY6iGSEia9hau0GlcPiVEx/Emd0T8L3rB6SXz2H0w
Hdpdq3bR0HNeDL5D9FvGk0OfRSQWdqYEkCMrKyI0moPphpcZWX9BAQIh6EQHgLcN
dSa0Qms5ucypEs/ibN3scXv/XLYoGSksmqDZSai16mfe/PEunTRE2VQdFhohfXIB
rPG2pa+f0TwEQHRmGe2MrScfCRufXbrWT8lK5NPizmOdTSGUjyHErzJIJKfNnNp8
IlZYNrF4uDue1i47TRPFiliI2SzpetkoFtBGdhO79COYwAH82wvojDtmZfARnc64
bYZlDeTP72VFJMbIapdlys0+hZCVb1Nmot+cYOJpLpIDUfdJKbZ+E7GcX+p7iuvu
/I6xCsZNwU/KFr8Jdj5vEM5hvWbLU3VlnVwwMIiS/35SmFnRCqwyPhByZ70nw2ky
VXmS4ObBhDo/IfEMVc335vBjocy85I/juEeTiS4sDkSkg+bi48HWLZOb87EyviRn
gappiqh4tvuFGX0QVrKq413TVBbKEZbOK39snpKVJkTjkfcxNvGLUJATCR8/oKBt
2u3dKBaJ9a02L+gmuJKgfnDBF73+DJAw5jYAn0Er439Q28DwlHseSBkFQxCcJikx
igdF+zepATJhdCxme58qzinjLP9KZX/RQU95ssD9wkNI42p3MdmwgXkp7O+QEfU9
7TPrT4a6/XKokUAnBj0kzw3bJ3E+KKgxlVC3DBBVWY39t0xGnjrUSS8QhpqIfA82
O7Cfj8pjX+MFwR+IkWQc2We4fTc1OPpTpBPypxz0gtl96bGUKRUd4JERPybK5ZcW
DTL3TTtfpqYlIq5aiMDzlC1Vqsjq6XYcautmGmOfBmOp7Kz84vC/6i6x2uRRZJPw
YurEjos/dc9VaeRKCBix1i7GzYjw9lgYpdfVz28UOBx7qgQz7Mo8zcuLZIf78wZq
DxslM2Xx4uz5VC6tHnXRzl8ZrkYiW9aY+lWzzKKbnV3wb0cutN/qovSvSxqS/y/N
KTDJRL1vCq3Ncwmt4GrfpDHrzWnbKNN6aobGy5Vfy6kq74WeuwaBRlZ6t7dFnBNk
Sv3p3ouq5Ulf9chp5LcVRkg7kcW5FCopeKm/QpIdsEM5wEsb4chT/cD9q/4+URtV
E7oTRi8KGqCCg0gRJq7SDsEUPBdLTuuGYPRbyRgHSsPVbby9iXxryljVVZ0BwV9o
WdVWt1g1DGLLh8AAhLBCvqCU19jOPjRoIqkvDeaKQYUdJe8Ze0iHVz9JksPXdJxA
oGyu8ZN99iZ8BRD2JK2i3z5Yx6aJGqIMWK4DZl9NZAJQMeobgHpDGWUXiinYochZ
WPxFgz70l4DAF1l3L421+HS+p5CYpZKxNsBqsMxKcrUMcFlT4NAE+0aEq7j1/3SE
5DeKMhxhvoiUrX/9HhtilaJP4QOuyQqnDFHZzEexP9SH7Fa+OaH/WCt/aI2FEAeD
CrCVd0tqxyvlaJiZZMGz9tg+Sa9hm7IYlf+K+xt/6jhKDvamdr4iCrGqjx/FVPI5
jvkHS0NidJG98/hyA+6aM0282X7r4l6SEFSO7WdI5hwXNeHCA+HJEKkq8ulLPxLh
Ekr20gb5mUpNC/N4XlYVst/DgAoALym6NSPpJfifk2D6zxhTfj0JnjaD6oXLr5FL
RUO3xUByDsh2qDw4cXz63q+NS+x3+T2IOsEWMyhgEE1UatDSs9PMm7UY6Pp8XI1T
HfLvRip+xfKsZSbWq8imAkLegmSHwCpE0rBHXxwJA7GxjfIfQmsaKpHE//XdLACH
QIW975VxuFsIVRnfgJkTF5YeRwl7VLHlKzn5ApBSSD8lXW8Idgz6LETOq+QCE1mC
jEjLGEua17AhmdJA0rI1pwHbrC1ysm0hff8VjeTxJefYqGaZnC4+pQkZH7LG0AN/
tJkEfJ6jVRGy6xjKP4PiQIaBXFxcn+5wrt6LUXJbX5pYjW3RBwBw23Hhg1goqaM0
mDq+kRA9hPmFitE0XJ6AHG8OBViK8NZuseBsgrqTBQv0JdKp/Hm+mlYk9wdTr9vF
V8zr8/ifXet9vPnL8fV2y7WNe4PaHXmQriJvD60uPZBAAX/ICudEKVGnjzzkRpzD
Zklb3tDboaR46ecZNdhbroi2Lie4VR+Bcsnir2kjnRZIsbB7gK3EYPCIi6ap0egc
Tgbq5toPSvICiNS0BR15lGI44GdXOgnpS+cPZUPztNGKj1fD9Cfvl6n5/SrgHwzZ
EG3VQhMsmjShZ9lyOb5reEiAMjZFlPXCt8FjHeh078vcCXtlKNY3MEvJXvwIZMhA
/5LdYtDEEvJQrbnN+zAlNaa9kaPgt9aLp44Y4ObFJxI/0Tky7eLr+UcwDLoZx6iM
y+oSwRLK8Ak9sQ67zfVzoBw60RnjosuUCmfQMNAlMNbII/bO/cvz3bx1T7bLwn4o
IVbspMpXEiccTPRm7/AUfvjibQr8wom2kaK99MBG3//4yi5p4XQDDMFNrRKWO2JU
hANm/Pz9EYg3BYswLSxDeXj2DaK1SUDXM2Bkf5Wan8PvEn5FQmi/yRE8LDy3dMlC
MiIveDb13CgpiZDJhDPxM5v+ftau+hV59xsIE6I4oQ+ZE8WOgGlwAxQ2+wcWkOj+
Q9QDtrjGd060X0CDImGKLqYcqz20mD2lMcNunPqBrnKntpHEupF8Bn/KUQbGoe7+
+gKzfZoWDnUlaVo6Ki1s9Ng/h03KtWy1hU1NyTowk2ApFH0DKL589rypRsReX20B
BndoPzBPBDNdZ8H47tbKdC5MSj4LcYMk0GZJQjJmPbogop+XhSIngCvpmkblg94S
T/BAZnI7O5LlO6nWe0HpUEh+K/xhC5blydidaiopmAVPFzJ0N6HsT42alokukjZc
+2chOC+qE1eKyWZqXiJ3w1/aQqdt4IurT5ux6LLB6zAGe/Aer6IFyNlQZV0zv/5s
BjC4RjHxjqGt4JIcVwUEpkpUQ28qzHAmnQABYerj1xrnmENLHSR8CT1+xbIOZAdo
L1QjZKdlUevQV23keHiAGUB0wdmgKa9dy9taDmmK+uW5iKV7NB8cEQlChh/o2UHR
0IMhv3nZNFROZ4wFnTpFmKK/bjA+5GckqXBZHv+5m/FzFcOho3dGYUWi96XURL/v
ly8tE8QOTziurPPhSjNjIbg6Y7orrzM/+A4tswearLLplW0xPwQDaHWmjtgkoVbi
7mNbT+DcZnIyRO2AgvG7Ghp5lCZap/Ft901hDHDk6raZgDDmQaRai+zYeOLhF7xZ
gZR8QWTzHZfQb9CULPBVqeAb4GfO7yuhQ4T501hXdSkRK0DXFW+ZxWtUFfv0EJ6T
OlUapwkc4YhAw+m3QwrXGQcez4xKgjRR8tSzKIh/z9NnmOkw/t66kRxP941q9IL0
QIZRCqlcCNKgnwUVtGC7W1YYFVZAJ9z7B4ZPGeSuul75LeQN3p3YA7q4KYhJKRw8
wWo6rh81iVpuRaZYwv5eTtq8rlmOr2HWUTLv7LVJWk9sr3KcOlpgMj01hbmg9DEb
+GxsPNoc+f8zau8SabXDnaJKvlGsSldMgl5tvlYtMIpyoV45IMbJW/pGr1O9uSam
0IHuwMUtGwvOeEkmur1p1hEMOX+THCB1Vzq9NvANQ1Yjk7ad+oRF2WZ/NuIqy8l+
KWFcyYjQuD3l34efYnFg+1A4M8uU+7ags8OvgiETh5bwOPma5BL/Hb9vQTQOz66t
7RxyTfItdf+qDlrNTpu8eJrWX7EftjCbQVxxUugp8l0V/fRsUQV5kkU5LqCLkkzi
pycdZVfxDZTZxUpnaUFb6Wsho9RZUkBOdfTWuN8IrqvdndQXm4++DAcJMu/ThFjH
X+/0oP5Z5KK6rDRBUFvTQLKIBTkW7ZOS/ck9kh7KSovZkTB2jKph49soYPV6EPOe
LquVJn5PeIlml2+NHOThidAEK9ng+2AQp0Nlgt430O6nWsiJ4SZ7VLCW7OQJ+3S2
QXBImakqIQ4dK3qGVZZpjLv17B/yXtr9bZCH0GpFQMnNowTebyBZeFq4ftFl0rDT
snC/IViYCBPKZ3m24MAiZCN6jMlMzoMXF4iocC2iF06EnWsAaxJD19gayUfzjsWs
z+6IwzHXOYqUvVt8ycxeM/i3WtaWFMR4zZshffZushOgMTXn/aqp8mPRFwENRAOQ
QOyCF/jw+ILCKjdaRJtpeG2qqNfe+E3lvtprUTutXbtfLWTKhxObn5kJVx0ESYeF
GJOJMeNIZ/fGWqDT5kCrBaf4DcARQVB83BV3LXJ4ZAmt1rwcmRh306q4xTKBNc6O
j8Hfk+dM5p+RKtC7MUGLNeD6R4FE7WHpkFFcJMPIwhnI/xfrBGjIq4CI+7xpFHQY
akxmlQ+3FNHWBzBckgQQEJra5cUv2Zk4aPqXQBkRbQgq0HDG/boPT0DGS41LM/R1
+ATEFiC1rL42naMvqktFdQZLOfBJzxAX8jjFSPOaJMZdw0DsV4YYhRCrvM85LLzq
xq2EWcclgUIxB1+b5VvToU7X0vX2JZcuF4qATGE1Y704X9I/CY5fBE63yp+lmyle
A3qKZZq+hftnNJoP8Vk1YrpLFzs7FYLkdp+A29HHL6kwKTbfRCeZdCW2HbCGm1aG
LdvZL3+CCMQB4nPOHZEjWb3+D7EmeaMyfoXQyukvMqx91wADVCeRiHQBMjWRCRNa
W5dK3koejfZjk6+SOvya+8GKtMYcTmi8JLB2AgIvggExQP83l0197yXL62SzB1AP
XbMGvaZZMJWFW7Aybh4iJ32SlO+LB3mK86GyNfUOJsspEs516BA5bUvUgzP2j3ID
C3iZBHJ2ITI8XMdmBFNYE7LNcqofktYu/nX7XeP47A0Jbz9srp4TyeG+6fhdu50U
x4vsdbhQcIQQ60DOkNtoyu1Xw580L9WjUPb4lRla9B+JUw7YWhUPGvHH/iUYcigT
02S+SdgjkuZJY4yCAMoRmeL1LXw5RgtFgfbj/FtXF8MOQrAbwmDFcbs/7JrwdF5L
KfiJUa7bMV8VJo4/60ioEe1aol0omrcQe+Ase1UJ7t3cH9/rRmzZ1vqU7K2LjLZZ
sUdQwLlg06xjNmXFGLaHG0u6AZS3Y7YOLu+DDbJkKHEo2BNsx9OwmuZgdGG9s/62
AadI1UvGFAztXVJwfLC5qaA+hr2t0HS1x00zPj2BRqsg0kmwGKQKXH2mKnFzyIjd
TQShavaIcjABimlAX48MH8f8erev+dY9iCdwjqlUGI1kKi2yq9xg6LtScV66fXzm
08JOO+R/rmTd/P9xGCQlRlsAxrg6B7Fv/db1kOO0NNySXIYvvkyU6NrGlvWhiDZ2
r/q6gyMDBAdOUYmbpofD5JvYupl2YXXvtQJCQ3OHjamBtaFDTuboZaInBJPJcz9Q
vuvaW/hbVk6yO9xsccD155LD2smHPzZPCndrQq4+T4h6gGfl25N5US5TyIIyMJy3
tD8POCorywrvk0wpwzAN46MOvScahSQaU7V5c/Gwf8pW3HM9IPQK1u9uvCpmrPcX
s+r+XviN/hhbcCrgszp2phTGOuUUQ/7ygF+ks+gDMrTEWPgWk+TBUGoSKN/ohRDr
eP1HeUneSdGmJ60PFfbPfgAEpgubSW+N3U+mtroeOsN/aASMyPoYh0K13FWrLHJ1
qTrioFVa6A5HSfGPTV2X5OkNeLHZSGrf9JyBLYp7LG/Y5/pDq54g2JxFDXG8sSce
9n2MDqrmqRI7JXElXHzzG0X9sDUXAup1B9vtMnocAWShP+4ubJw719TTgkp0TAeX
29DFt32MIGMAtZ67vuosNBp/ZH6B8+OsZdRkOINnJZu9acA/QcHgYaTgMOD+KRsQ
GKUUPeVyIegvgQ1Rb+luovQ6rPnJseQ1eAMsZpCe5yPrDf8uI70MSg2DYBghYeSK
GWnb6PWW5+o+no+hnhKCnF33vzLJHuitk9Qeq6HCW7SbG1dwrJS8GdQDukv0NbN+
6Xb1oDNK5czF5X6o31Ff0ev7+Un05apa94KIoqlSMCJSOQ32HmU7XXA9xcdcBnv5
ONjzHmLvlhr+ncdcKPNlqqtvxKg1VoWuJS4PmGG7daR2Eoiz/rOYhHxctvsXhwy4
LER4myzNgiC+gANdL46CXr4UGg4cfl4/QqjM+7Exb5kD3IjvhctqkL3Qylufi4YI
vgJ4ssib/wVhARN1MlTK2eKpFSQ1u80Wk5nafDi5qy/tzEbf0NEYcxN6X5Rgdizz
qg2v4wAqDxbPZY1kAjMSc8axF6YIKW/1o2LT710d6lq0+4BYyD0Nb+k+YX4NTJ7b
JT94dr+UnZRGp9jOi1hlXer68rNYJXL1QZIoAo3kEqAPm6QQeZorFl5JT/tzIP60
0OyGRD3coiguxOsRqwthVlsnfA2+Hsws+4Uy2G/TmuWapyjHEpRTykRbibQ0lbTw
NwiCSUyxEYocJs3yJdV8L1hTrEKqytmng4NwpzjHUpb/IA3u5kSUCyh2ewjcwiw9
aOl4BNL15qJ2iZdcN8cAP6u1SxUhInIO8wrdoEhd9rakSGO/l2P6rIrNFOCgvWr/
OHJ0p8oIMLrEsaSEwVan2K61dHJU603ZJAKOJbaPoNV7k2SMyxAXlIlahHObzc8O
iR0KjG61rzq8MaNa151uXQZwOcU9MMYjvIvn85mcgJe/cxJei4FnqW/8uKblTEz5
fOF59Ywea7dzK68l6OiVSUwZNpMnsTnQoDbxb6hz/7qJ+QvBqS6xX+STPla1Wzu3
2SsArLucNgSGSI6vdbz1KL+SyUfXHKlCwDEDiLtmPdBU3jffTZHWHG1/FrZxqpqI
anw6ElgAKNXfMzOLxWRsCQgzb8ghTHn2F+qAs2br7RLufGZbMrCY5pSjtPqAJ92u
NsX6elkNjWdDNo1N1SPscQ==
`pragma protect end_protected
