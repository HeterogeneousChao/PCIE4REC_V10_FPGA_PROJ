// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:25 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sBvf97LT8xbGgcZtWJcZOTi2Wja3CP1/sdjh6ftaW4vr1GpTyf5N87eHZ313nSrV
ED90iPccZPLkSQxIvgMsVwN65KNfndbFxpUogYE7YQpaGOkTCmzfQPMkbdAYhFe5
jY+YjXFv370AuXXx3mm1TPRPJobKdpchdxELWvRJXF4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
6Jph014pkGv46vL/OZ7U+htDMLAjT+uJdOFZDUWxtUGZqz1+WUDTgZ1cUCUurEfa
49SNPQ4eHK1N/WoaW3yrWQSYY4ZBJcvjlVe1lQBh5pbBa5vJtFCwTbcX9a/5ssyg
YAcm9HMd5wWncWyE034q6mB7FTeK8HQzhNaTIM71shn0v24gTWsLDfpt8g8VJfc9
rgZRfqtDu3y1tGfyd2I+qiBTvNeVwZZccUTk6STo1KjleqsdAC1JQve2Ax3UsrjK
nfKMqQGvw//EPi+M4c21HbJPePoCAGEKXMSB774qZb10PIo/aKR3mhkid3qVGbG3
Q0zd5PEiZk3Hmw/2NBRpNV9vTcOv3OJbgAy5dMMDwcKnCB8dou/H1MxLMfFG+QJ0
15PMEMuLK1QeZviMbvhbJlnOzJQiPUhjAj/ZDA3EI3kg4P4lh94RkAfFlQOujqbO
RnnN6cnhfaV0xWVcEerBDOXlBAOfOC56EfPy2I7uTaDDsWYTdfL/wUTeWo1S2/zn
4PB4BpRJ9oVrb2Kf+JWDq5kLk9sEQN81BMWQayFIPpcAJqtz4yWrGasSXBQuoASt
NuN6Ckbz1cHafpWvmLb0gNY5bpHeU7Jzq+jlCAVQdgEo/M7uG1eRULUx2lxALvYk
pudkssnFi9LkFoljpRvAD0sMMgQhOT8gwT2kbDXK5rUlbRfTJO9Gaa8+12A/jePt
bJr+YPsHiqhsnNnOoTRrGmuWwP/WWBl9pAxTKZ7OHK4sARyGpdeK2bLvigc/g3mF
crEOQ6QqWVjUOG39XFRDNDp349Gdr1b2thHM2xg5QWQr0/WcX4v9WJrVPe1MJRiY
3YCQrjbgL3g68lER2TsW2e1Dy7nyUHXEzx7p/dZqbWpM14D9bXa2UJJ3h/01kva2
AfbcGKlE4SjZ2gEM5xHIEh7g19fPB3l/Cur8PFV+hokEWHLscYqwe6gbGFsHaokW
E57xrJSd7hFH4kCwUhTL7jnT1/gXWf4RXkHto9NRKqGcshS4iP2FnOiGoE3Rrkzy
TSdYQj0snudJyUl1++nckRnkL1DPq3sgd4hCddQs/r7REPYtx3jDwGcQgLa/9Pbd
2Tl1/Afc6L0te72rOtDZepEyKhgrhlooYVE6SYPIBgOfl//ip7YKwtBaKzLvtWSG
bNZMuQbxBsLqABHKhuHHj8anlLmUUDmzM2FIB90g0y1tTkFGN/GvPF4YX02PrLHv
YDnbq12ZzIcgLxHKzISemhk4BLKNR3zl3Df01sjh98lH48lvoFmNyj7d+m0a7TjB
zXtOouMTwLZh3t+KidDItbFdB2Jf/dOK4Eu0aYscu377WCXupf/2t679OXaGWzeF
Ocz8EHqLcC11xaJYaaR4CZVhRKdRLWls8rBU/rasNtFTcNUnNThmHGte4Id7vQyG
2LzRWOpnX7i5SEoPIdQKmL4ZsNLHwlI6Xep7kngTIgTlw2N0vMznxBmI6cYV0/+Q
vQ3hz7I8NvPTFxBxC8P/NiOAZOoZULiWijWaHX7KG0pYrhubnwhEOIPlnY3l2WW0
0zY3VLR9VqUGP1oURWZyCYFO4NbT+7oBzU3nHEaqBxeJDdRGmAkeqDgGowoSoaPk
WiQ6fxfEgZzLaT/TpNm97649VNrtrPT7PCxNbD8pOmmjh55psKKGCHWWD83i+84F
ZuvtYn0MO2aFlzKxAsAGDtlr6Q9c82aTgc5EbxbvniojlGWUzknww3bJ5XpHb7Cm
OjhDnWFpvNAQq87Qf+Uyd7Ds43Z/Wh4S47vnv5DQDVe8hcRgtLItyj99lh3X5JZ5
NrEFs4LSx/k939zp0UB4yPpfPsjlx5Dg5jJnzTxthQ6WYGurI7V3YGPc+PPJoTeT
UURMAgt6s9IW6QDWwBagaR/JKW5n4RtersvlPyn7nYsXt1bI/1XGVN5oXg+rm+Mz
GMUp8xOEc7zUiwx5+6f1oRNyD4zue6+mEwZ6j8QJcA51f5UF/Jv6GdqWLqtTCqih
QgPxxLllduTfTAT2vSWyjuOmqFTpEuGE6CsMN3O8MQxUz+D+5Xkau6dvMgm8WYuc
TJJFbHpm6tJL6Hdgu3RPVI+/i8wD+K++tJp20mkAHheCiLHN9m3PMQtqvq6CThMW
VamwCFpYff/bSBUQqMxU2jpHBuuOXWSzQsonqndsSS4n24icqiQOGYkuxho6UOGg
DC6CwAITOY9pZm/QjjBaVxf68eh2dnxCc0UIQfqnrPamuwMuHyPeITx38v8g4PcW
02hna10NQCsO6+lT5OdMT0qfy0qkxtSNcXyp7DuhJHgpXWGn1C/C4xHoN1E5zzft
SCuaEGSsf3kYIBRdqX0eWARVfnRQy/xNoSvXiDcxughChUO/1HUak5hw7cV3Vi0c
jqrzpUHyH9ek8rtMCID1nt5qAq8qxZmmjzgM3r4ecDFrw290RAQX5NnBHbrSxlGc
PnQpHt8XRUgL6yb9kXc/1ZpoZ4JQJxEro1Cx9ZyUR6tdHUlmqiajIo3+WEh/aPAj
QVS+feAeRJAFx6uPcH0slqcqI7o8SyPzmL0pSM/XddvzxYsCUcpO4cJWd0mz4Kkg
TTNgDWifCh8Uj5VQF9U99wxckeBDkE941axFGdRVOyzTOcpWj3dvLbtOitBzY7QQ
7ybx5pvzGZXFdanhpFusBcaO8aGjaOyPL5HnggOE4tjKC4wp5s6ulVO0jmgB7P5l
y9c8q9mXbSp7dqm1P1G92vRsEI65tqkLVWIRif9+W4kgNgOobtWOw5jsVCDYJi5R
WDK3F/fhXqG2PiKiU2r84l6PmahAh/hfjYDoRWEVlwPifYXzfIZ1CppBqnb3eR/r
xDH6A8XOkMfwwNzM9SDsvvc7JsCU5cHOaqrihmbFFPhAUHD+aDUf4q6hlFeJ6lkx
vm5A0c8V7Q7hXS1nYGglNgyXi5tphf+mqUGm/5d+L3pzin8vR4NQ/J8g3gn6mvmX
Bc08BXZ1UlTjlQHQ+bxos2n4ryYbgrFD6+l4anP5cxkx/uKTRUKwF21UQD2O1hWI
qlS5tUoDQ38IS8OCeNaUzmoQa0iZrG5Lne0527MsfVp5x9n28Ll6VxbTeYdgF+Jd
q9FalVxpccppPJ6GQs7qoEfGOoWop8UDfy/gT+7t1TdseG5GMCSE5kUGi84Snqnu
aL9A6hTUebcG8OwTkSe2kIdUZujf7X43v2vFzw4c+siFMJ27Lz+4geHLNoUpQ6qq
XF5uulX9+ccuDmxlHdmoj2ZpGUVYwPe73Z/VLA7OLtPRh7F5Mz+tVu3E6kVrb+Ma
mUFPYTrjpsLTNeZC70Uiy40WPE7SyJdMG/a8pz5AWKGD72ZehxT8RZ54kkuFYEdN
GRXMlAr4voYAT+Qa0weqw3WZbQmJgDijutD0AGgwK6j+nHKE26n4eupfE7dfzjF7
wHQt1M5MMCwpjJTYFf9Pc/q+OctMd/IvBOns/Fa6CXsET1+6IUOznsE0dStVtcqg
Ehfdo2JCjKuBmyI17UguYDUf5v15Dq+lYYJfvx5hDnmKCqs6lXzVpmFAM/AGEZTu
m2+reO8qhhHeQb0KyqpPU48oqyu+EPD/exvOqxL1QFcdOnVlqRJkhUhO3L7HlGHT
IDOxvW3Ip/lB/jax3uktnQmnWsq49TZdbkys0qQNw2utmlYvDdGUyv7s4Ent9Rz5
2OZB7e1g86uo481gMLRKZGjJkBurp1yTiKNyMvp/RV2P6KYdGCbELX8HEjdPS204
jfbexFBn+G6geAYvF3G1pBJuz2OmmiVAZBT6al1FxiP/FI96f1mGM+YYD8wY+vMo
5h1iDQ3iMmb4kWwtLLQPqkKnl6NUrnQcVn8zJuCjV7tfOZv9h+8BGfCYUd1ntPsJ
/SQjV9nAHK9oclPP11G3VOBYNJ53a0hg/UbobCCSFguniwqNOC1+6qWpB3Ysw4jL
MV7ujJMZeUETUla0NqdbltAZcRFiGiOyeEpcgjTqc2h+1+pTK2pPLh0Tzcg9yBC0
VNi0zwjJNcICAJ44RhGPA6/MrKZlmR1Dk7tB795oQtgDKzIXhZck6zW62TfK05lX
C+mRhiANm8VMwZszPO+kuGNm/VTKaakpYM4uOMovlotsz0g/fdj9G3YgWKLOLLu3
6UTYgKolnHaLgRX6+2H4t0F9L024K/KYMMQe8qpo4bH55kwfIWzNCw5Yv7png++8
RlJF+5OQaKSvOg2HO0mMLsk8Wq6sMhu6J8kkbq3+KIvyzfBcsi3rQMP5ZUiFdSrd
fM+VEc44F3On+IyRsV9Wn/uMbKp0QSYefm3t04NyO9bVr5+evqymZcRVPqcY85RR
V/GP6k2FimxXDjv1pvqla+Al4Nm2bsME0Kj8LBKdazQS+h6sC0ye6Tx1ZGkKUMOe
JScoCm500oA+C1qTVKutR3HlAlO7xdsIuaLgGrah1lLuCjQjXs5kOqRiiypUg5jS
vVtwOZAwdjd/mFTF/resk/sIg0Gs/RQSJ6VouNWU3SGXP1ajHTjS0ImhaJNtg1wn
FvYelyKwNttR8SIExAT4bkT/EYxTCLCgp06x8we5WdASx2xb7bDUX5SgtrogkS2W
4u5DA6NcVK866vhTM6nwCOG7l642JT7toNOLGhUhBIn6BOVXQ7TXAUW8kJzwKPCN
YtMLQm18bsuDJC/3AHzlW+uBKFhaIC5w9IVcmrddczNNqTeG/QB685ujIk1IsKhQ
ZsJghwKm17DT3PwRCH4n4crjh2+Xp7tWVzonhmudK13UKKSpbPOnGTfO54Q1OyHS
OyAyc+fBGxg4DVbSX43smPCkjtDXk7tWdZHXEuE2+hgnC9siL9RoFMy+babq/VhT
sB5M9RcNxjXheG4PPv/LoK/XD5eTagfsFWsfhhn2HHikKhpnPBpf6KmeHPZWyRhZ
BGo5bIaaek9OWtMyBOO+4rlEQ4iW3yygQyFpyWI9lFoArWgbgm0ONM7YFRnYb5Kd
LFnqSs5rSyf6/3hUH5aEb9iSh/V8cYK0GGrS6+F2fwa5WtF5AEePAxOAuMuOt1yn
wK7S8bbVOWZEAMxec36DVtHYOQZuGagA0kTb2Fb+4mA1Ccd5tkSpUUlNSGL4YTTb
SnxYSL0O82L4jF+c7I7JShj92BQuIZlKcicVOPnDDhbnKTM1l7EOQSw8QFt+cwD+
xXUe6hwh/992p6CD+YLP3vsr6mdV9P37AbC4TyEAKitTbe8CwHRGpIgkDSJSlDNR
xGz9om97LEZbCeIfEb8s8AxtVB1X2rG3lqfbT09/AVLg5qN97SkatSnvXsP0Kn6W
FG9wNZFXgobCUJWV5RV//2KHGFYlKxThweb6N+v+9rjlgbUIVGyu/Rx861z7Eu2h
+tuH+4q4FBiZFORcmSvZbKuSlS7yUErLMcylzs9xYpU7JkDYROlWHozKxP5Sl6aZ
eS3BBwoD0u2xiSJ7EI3BCt4afDRrRn+my1u8bx7Raa1FO/4tG6Dwpov7/SKv8z9i
3BvXGP5zqvyGNGjTc8M4bHs8X/objacQnP0EAKNOcSTSu9Qws42N1LiKcksMbdLP
CTCQ6ZY6oiRrIFo2dFmxzMG130LqGtfOivZ6woA0D9iJQt1Zo4jO9O3COMLkvD3/
zsYhcvQTlk65Dm5Ehv6tBkkvC32U/JREK68MJZWbc2j6qb5dkw5oXcKUafu0Fspe
Q8Hte1VNoeD66IPXfdqGEvsm+bSBI+jXbX7jFLPI9Du4fNywj3kMXL1HLVM42BZz
Ds4sbZ8UeeH73FyM/BP+ryBSGszUiEogFBi7ZBEhR9oYn7nQdq0W/PQzSoXGNX7R
59UVReFiA/PQ/ot9Xtvo1+N6smXqJDKCi9+dyUfgS4Fgg6jmKuRj4LxGQ0uNiYVR
4A9abmI6j9fqjM9KVocmyt4w1Ycwj9p9qsAKIw3/VYgu2XqthPJhJKEPNDloMiwm
1JPNLrpf+7SScRr+VtNhtZfTDi9e473wSGt2SU7Zl9iTMR488fYtp6SqZjOHn5/J
itaA/6bVaMA5IPZqrezCARKq/nEuyk0uqwTo/13hadgfOGeWGML6aYt90lLOOb85
mAKlCR2NhQVFspxx5mDEJJarUlP0tqIdLpnOPgDDsrcsuVYSXegzpYFVM6Shznu8
0mdvmp5yiIKgGXl0keu6N1xn/0jmfdkX1XKihToBydjyGArN588Scfk5SUivQYpA
kB/QbSDesJRr1QYKJq48AJ0upmP2U6r0xG3C3lyrb9/+ebVDjgL7eKiDizgpLW+Y
WkFAyr7iMIeQghrx+uUyXJwScldbIWKuXR8YN30UFfLhXVsWPfXFYTMmnCsxa+pp
B4ktfrPRQwTd1nC8wGzjEEyQ1TP3+Q6z8gqgib597ZhROrTGhbLFscbAW6Ccu4th
C51/hmogMO3bpfHo11L/BDPYohM7X76AmxkPIgqA0QLN68EEE7UwZ2PfjVyD4IH4
xzcKoDFdwqS5bOx8bgfepWfhiC3FhXGRaLP4Wq4nyZE7Z1/AoDOZZIE1cCezdYNT
ILJjyTQ7JiSu0vlnz0qrrmfusCoTfLmjX7FcLmkxFocjjWMHga3vIBGk8dcn9Z/w
oEc1rtodlz2DjcsDvhuRE8IIjhXWe02r610X4n7GUkP3aNhrVUqzeqtOh3N5QsjB
gTvouo4WlrfwULEZvV2ajd5yS0Jcbxb64APkUGi/wpUNgWplXR/+7YmsbBERQbnM
na41XNKH4aoY+s6c7DWGy8KO76Wj8bfsVhZaS+2Y/AFJiiP7Arj7lWAYm1/PztBN
1XEmlgc1E78z9okHWTBf1ApJ6Ih8zCjRuyhCPPk9mP4lw3r4G9JqP2Kt4xwLplWR
u5chKsEEfFq5bL8Xo9/byTvjrab++pw5LycAgsL8QMmV1SiO5LsH7JGNg7ZI8X1C
buYxpq4Jmhh2u3dSmsp8a6p/5ngh01gupTLZvifKbkjMt5i3QOGoGlItkvKsJx2R
3F2X76UGS2eL8didPyGD5zjGW/rVBcOcfQtrmBr3DLtC2L17F1nuW1rDzMJ8vxah
QZGkRH29CH2aI1xjgKYvXEtiiM1P+FAQjGNI1zLtQSzKQqP0kvHHfbdbQY5PLn8o
JCjpkAvwTICd2932HXf+BcD8lH9KAcK89tGuv11nlUsGGT7Bau33gjwEXiUWqB2h
lMofkIpCy9nR9c1/OkA7kwy3guQvMs8tpot/r1nRiROIDh/PluDx/XVgGJZvDlrB
nYIxGljAQmR+dEov8QgFmCT+nSkpD6DzP94lQAdJ5unwvxgI0V3DFO7C02znYKd4
8sh18UU366/PyertirnXuiHpDS0VSLQcDMZxGXhq80YeRuAiTPWrlT1bltBGS+kt
McZP4OcwkplH5Vv1V43vCpv/cqHT6UsTPfZIUX22llenvjcbBsMAGUFluqzspxwj
ZGXlaEUrTkocbQ4Juks7XNLtI0z92NQpcshk/WKbaASANS6NxsTrB9lvcudLK2VA
DINn2HC1qGlRSi0ZQH0FQN8mGOEXwamWi5nz6tyxVDU=
`pragma protect end_protected
