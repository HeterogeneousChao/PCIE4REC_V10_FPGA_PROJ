// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:19 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RfexSJydCu/4Zr8R22SauRsQ7NKZm14Tzq58cIVjNpVvpIRYfSBWyPHekEOlDCNR
dRF3VJOSm3I/vm2W9Q+h3tnTc/yhioHFNaoeDFo1+UCXfafH2UTPy/38wIj60U8t
80lfrW4+dOrEKmh255S6MB7cbYgEvTBXH5Y5U70gwwI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7232)
wFGLdGWrR+WJiUGRbovoPf0hnDi4oMo9T2VfveCX1+ZaNFgeZcuC21r9Nz0r6Hx+
4IIQTyNugkVV/Js/1bKZK7J8HsLMNanYBBQwWzthtw0TFu3JGSmkFn1sFoxKYGiR
OR3ko4alOuxy+TjmZUJPoRjlSpsGEqG39LEJ8m+CbZ7ItpFk6LqVYfa9iQqX9pak
Fg5qci+U0jh6seiTXt+V+LqaswU3WrO6I0QNduA38aNJ7t7rs24AbL9ZmKVyWOyh
igYUBUVUJwo7A1zIsattlK0Bbzv8Cms0BfOL7FSoCfWostfu+7s1vIHxBqvvmxVg
y1H99pX/7s957JKvK7X0rNCUIg92IKAagubVtxoK+SdhITm9gp8Ld9oYnTSkazmR
eRby+7nCoLStMQfuxW73eO1AoJQXRlkM0DqIesYvXwGYXklYOMhBur0n8HR5mvRH
xAbgoTqw1DRADq424YuWG0cVcNDiy6v3w4xSU/hqFZD0ezHjJ6GxOXbymlUAxA3D
g6lJUz79Ht8sT9VGHDtvN692DS2kfbvvxneeDw2NxlCKBAG9MjZvNX2IyjCLs9hF
lI0lGGsvsSY/Pq+3ProGNKNG3tAq4U2kDuzPa3mu6YeyOFEGxhSc94tsfalQG8qk
+U93ib2aKvEHLZmttRN5Y1HESYuqCuy1k7nNIexlDDnWAbvwcd9Y7uE0K1mJjlTJ
y+WpI9TxqJrZyWJTh/Yb7nDexXn9Z+Gi7FWg/IWgOEM53skf2DKy9hJVZ5Ix7T8j
s6zQRxOyu+LruVPRIPIxPGzAFzIAXvbk7AjbJiFFPWWH+MOfVRSl1Ujye4si0KMH
gdMxjZXQb27ThfhWRvJBk1QSZZoLU29MoCMrtaqfgn8Z/y7es+zaNwd9vhpvL+6R
vakkC1sFXls7qBWPal6sTl7BS6uWkBcotsnlR42GjhF1kc/cnFFGrEO3h/DDP0bx
taPTHulu1xQWgrcxgbGPcsbRZTBYDgAodXl2Cvq15gTYhgqEwPUe01uDiDx3TTK0
aDIviQAhaC4gF5jaz3rDFvn82TK2bl4Cnw/IVPcgtJOiAnuHiounw6Bd9MYhKeG5
Myy4/vTdxF3HGEB4KIg7XUyg6omvzJHWLwTQ7fa9j58gpJNiTltmOklMMA2hsvjx
RAWDrPWDlO7ksZtmDV2Hyia2GZFoJrCUjhlOkUF7eEWf2/K2+ZOI5Ga2WpOodB1x
LB34BeVMnX8ZyZirZXZ7VG4eOREt3bcbEiGzncxOu7loyiTxmU5bjXeqSZyfGvwo
9Sw79HS+Pfg2/zVrHNYzMG3LlHcGC57edvqEhQlrMOMlSOcefqZTW1Y1C4BUdieV
wjr6THM21kFz/CKOr+4EncuC/WIRjNScNOt8OjXdunlvZ6JWzoZggI1eNqEghjsN
w45UM2fHz7Ls1L5bEsC9/xZ9JaRCiWXCLMTmN4H1r/wzG8OTJ/M6n42t+EJLyX9z
SOE/HfShLx8hFdpDiM6ZD5iX+tKMQuh3G8I8A2nDAPiB1ZFs5P9wU26l1fI11Dqy
fYkJThiHGr5O6Epz6xddFUwGgGoPGkwVhAoQ7Vw8AG0MWaDH8DQJ+ZJAUQzS4gdI
8hzact6q+8UTsZelP+ksgVnSoi+673vy/a2F670WCzI6e0TPMMuMbjz0YCQUxWQw
Hmf0KvdCh5zZOBSp50ZZHX5GcGORBGu4/ZWwimxTzPa1Ww2vjOVtyl2kKF0ovPoB
ec+AXb6+qV7/BYNBpHOvNW8RcpDVqJ+nXnvn3Tw3Ym/kFdSWj8hR5S7FgJBht1s1
PcPBP0zrsAxz7Qe3Y6tzNowkxfZXRY+DGyydDBWAXWPhwQ6/wXb4afuw0bfzJGcS
0pKAt5ZbRj97Cob2eUwguUYGkpk80o8uLaCtwp9XJrip2mmRtqZTMoU4C0UBJQNJ
IkbY91+Hq/BBOrAwnO3TfgJzSRZXjm6O/AjWu5QuybuTaJ3/JEgoh7Lj8Dx9dcpE
Apcoh0+SMJnAFM9f0YRj/6c0uwB+GDnjqQzLIKrV46ftzDWALAWk/0NwEBpwKTkz
ydEpS6U2VyhzxowBVL5kL5w5d1MJmAzFiRwAQSC1idHnlVgU6Q8eN3h8/vMmS3ZX
zEORIGOqpIxAZyqYWxMYREI8fVChkX8u1hY3sbkfRLMwR0yMHfSaIXVdM/NUPRr0
/aDXuBqOsr3zWkjcqEJAEE4tyzThRbQJzK2+pfdyI4m8abbEEkqUuEIXvHIM8JVI
rjvKyyAzG0m9N8I7NzlNJ/YKsyweo7X0/KozwoLICG1BP4RNhqfZ8XrBuWojG87b
X6ICO3QHegI7yB+FHi8HSv8n7TPNRlE9NHmu3fjP5n3zhJbMpkzBJEAjz0yJJEFQ
CXeHBvQLERE70fXoQrEMYIlOOqKaYxytpvolyfGyWF+svNH3L4bzc0nCpVzrRK8W
BedBlto1BaR1Vn2A67tT1coVOeXMVRoCoNiofc9FkosxftoRuukrEYMygGDg6UZZ
4bbZy2OCwpISPXr7Wo3diV4WdTKARAe/dsS4sJu8iBjVLlM/NjUJWnx7/Fy5mlPR
n+pimBZ4JOly6s1bGnC6+4NlDziBp8WPtZyvTRzJHEiIpk3znHAcFWsTQS2818tu
quvCXtkmHYZJZD0JnYZh7izyP+wrC/7C7b48hj2w1Aohm5jmnjYOpWbHLEfCyr3p
/Sy/3INo3jdQR/IPhp6Shz0xmvWbnxSwneS5V1a/XXWq0V+aM6zLsWZKrYZTeDXb
FNZodzi/EWaRsk/tJ6jmH3YGg7uVKYEfJlfA+5I2K1OQwOIbrql3g/R41ImpJzG1
v4EtKDZCQ4aiFDAXDFquqf224Qnd2wavEm+8yHxldTlwfdSSl1ewd1jDbB+SEo39
14GtXhRdnzNJkQ0ErLPDyld0yobk8PwTMorSsKXHfyt5qi2NufpzSZZ6zEZDq9d1
+Yu9wZIxS+V6HSj52S7rP+BKwDvdyyUDP+seou9gpE/p5h52VEkdmp1Q1wlJkYdZ
PyXlVOb6rRsynj4f5ekN8RWRKf4/MpfH8hufaoP4iALtrcakdFd4NI6Nfalj9MMf
faDUR6Il2Ctp2zOWV6e3xvPCI3YhInTjxdG/lxOMvbrJFcODYUisj1XLMlL4N9mv
jmqvjAcyKOBCs6J0eb9zIiifrEcsSswsNBG9cNsXPGNdW1Q2F+TpE0DOIATAsx/K
D6vLgZV5d+o72YcNSH/m3UaQWd6O0fRsLhjaiprp7Zz1bAiQhGqWN4Kyo21/ei7G
9tfyyLKAznv+UI3K2uAXEXnnJa1B05FAxNkk3C3H5UvQVh1aDo2zFiYyi2Nhzf36
zFo4JgGynXIl5YpAI2o+ZESLhB/CDUV2ty/wYgKutp9a37IA4Ai8Y5nekBCWXsyw
N5PgFiOXkfRiqAPPtBaM1Uw+KSAtYR6w7iwdQmv7SQhSuvAtiT9iDQnrGb8GBd/Z
PAa7AQ2iG9tgrFcvAfJRE8xX0Fvyrs5MZzYYoj7w/fm6c6EtEr+0HcW0sH3+KCcc
NHIREOKWR9zfeEm8DJOrM8h9K5ecIjH3CZag0fAEk0EDl4UgX1CnRviatPxicOm3
5aj1muw15WebhyrD26XTPHa2+8FpzggvjT6ILFdGYGGhMszhEbfLQhWdropJw2r6
zrfapUw79iiSStZGDByXQDjEgBNoxoO1W6koD6Fa2q8UNqPaF5TNfyKfcVpqE79X
N/gDD0yZxtdSvtSqibokQB3t+BOL3eknMtbiStUtayc9wIhO3eKnZvRuIq4pLQ1o
rZZm9REfLKbXnFew1aLSKQF+ETr+ofJ4VUSb8C74ICilWdjdgZZJAJQ/mljoOYLB
kTTokGHJMnYiPF/aPwXrX7lLFVcTonw+F9VlLfA2qMhrCY1Upft0o3AVbeU4WBp0
ecURrvmo6BKOwmB1MZPvwtXGkhJZNF7iryGOFGn55FoW1OCHhJ8Y8WNLGkgi+n5h
kHwf6cxDK7OXpWbQ2t67sM5qNrE8AlX1Swl67loGTEr25mn27r0B5cmJzJk6F+Ir
r0CiiDcjbgBTfsK9t3ymidrms+1lQdzBF5EuZiL7dzhs+xRZpJi5Um9yiufM/Nwg
hQIywDoLi+kGCz4GCWf49HwRvU5HN0rUVdonSONvZLgPs/MPx8OjOOkzvZCFPpk4
B6mfrdA0L90LSS5GK/IUVa8nAbEindyB41+qISyxcJupZZL9bEp0uN7atLmRmK1z
zFMZbmJ2d4aFtGf3O9f9WBoPIL2MN0v/iGtK8GoOZl7P83AGWKqHMz+jeSyI9Og/
yIs3XHDTVlr5ApfwyxLR87bhDOZZUHIIVD/gB0gPVwxC8iZmnpHgNRXk5UQ5fgSm
beStIQRbywL8h12nE0bdhgBaGvKguNkdGl67SMi/3b40FKM2P2vKW3LhkaBPNlNo
jJOlX3Y0fSYQkTLN5H0PxInCU+csj5GnyEPrAB1q9qBbLvv+j+i8cI12+j/Vg5ZC
gAZNg7LsO24lUqpRkOIGqShj0b69+350dQSESsxD//0EAvshbrsukZ89XPVgjIXC
g00ssw+GaSerqjyNTUUefaoZceQA/cFCJVvyZ7dVcC8pnvcdylicJk2eFdrNGSga
nbsOTgugwXyMH+sXTwj4UbNwtHNVrmQAjtn/+vWFy5vTL4i5tKAk5SG5PAeqv1tl
egpcrfKW2Jb51M2XKyxIPja4LS1SaBg7TbDS/A0x2sb8l88COZIJuOlUy06Yq3df
yrNO1cHMgJPiUJ+7IpExx7hWTjM1PZWb6ewtqT9Lv3DaCxfeUfZx1odvGhuMcFMq
ZXKZRDWMm55flv+t/48vH0HNaLQZjEPkMGUmX80HoEVUIFvvekaf2fCpy3bIC5Q5
ibk3GZ0vDrBM82KCIARl0Ytut57ezZyvWkz4TInInDu4EAeVp1Rozl9bpZCL4MIs
W56Qcdv4tjDq91weQux+Qq71Hs5JodDQBQ9noqLWBqcZqTUvDNsZTwjR6QMNG0z5
YtqzJiYpLS2Vv9yzIdVkr/HvixItjAa2RlepKNgs/ypsJ+OtDU5ffW9GmQ2ZVy/J
Ckh+8mlx77ST5YG9k8EAi+nfn+YfSkvAA0o3p0jGBdJSs+uxNAsvXbGW8Ap/7gHO
Vy9zft7U1+e5nt8re5ll8ulbi/D1gDlvWax01So50OmZbudVIZZwylzpqDsgAhbf
4J5/S+JGI/qqYmqphYxeWUCE4dvhC0weJyig4igoDfl5B4gSNvt5na+sf2S6Gkj2
Dv87h887q6eIeX+JKdYAHI0QKAz52aEsFUl9taZq028UhO+TH67mx9xixAanRyXf
ALCPNFqLwSksyl47Z6bERxJHZMJGWaTNzXNvNGR7jG3riom9BgmVNlrzqnsiJ2rL
p37Ps39Rcwg+v4exjKMn0K0Urv2caBvhlwMkvtjK2uzIKpbLWlKuV8aT8vR2uKVB
boYHdAFbJkzqHtxB71EXGmp/FZEFZClfz8YuvdAl3FbEFOMZSvXDv7ogmqWU37jj
3lgKToNpLm37PI//GCkYVaQr1BvD5GmBUFdGDAop5S45b8S9MeOoxntmFCK1AUPQ
7NRpSWFc4jrzB53cDlH6+/xV4AU2DpSNlNJ4g4Z/Be5ik8IOKBBwU3CMs1dOkFMP
u0DGwcNQpLjq6wYWhLkdZrrz0TcOIv8JqgUlehj4I5KhmvTkZEgFXZOQQWbj8l63
mb5l6yEr8nmg0EUmiL08L2BdfhthWhfN0fmlftssQWrLd9mwZfxKPuNqmE6ztn+6
3fVXbAL1MX8A1tax+PD7RPXudKMAo1nN/SOcf59Wo8EJN2h+PUtApcqFZPsAD+E+
3F5j4lSL9b8Lo12mAZXLm26vvK54g6nmPfziTBMrjMjgJHfL9+XAZ5Z9GzK3S1bz
Xg9D+9ihJEVRMZXMjS24tdwU8vALQU9vFCEOc5syh6MSwWJdsYdociy2N76DVgYx
ra7wXR9Isq6k56aUWqIg8CLHOrD0I0txoR0BbBh/wc3o6rS2gj9c33vtM7qq7QBH
e7QzA6EEk3j4kjiiuCS/yxXynUii9v0qeE7PPdwOvTWm6ZkV5CbbOAFNWtTPcF6i
49OVF5lKAnyHgjLqzKDwXNMYx7/GD1NnNGxik19BW3QXZGM6M/53AjdTqxSLwkVY
dIq3xq6jIBW64SOoAgrlnmOLSeTZ781CWp3h0O/kMLtQaeogCRCkYcZ67XTyjiXm
+tyH3obPp4b36a03KeYhHgUaaScwEP/dZMMjtBmbB1UA7iKN548nRIuqo0W3qHw4
NsJ8ixE/AggDLQDadKfEAL8sT4q6Bui6+BU3wqK1Ps8zr/8XBCSHGtSY3yvYhYiq
1zJ0/OFkr8MrWz0K9TMEDD+nSxM29Nj+hN8SpHneRtZJYzAJONVhbs4NF5AqdKo7
FhhGxcjYxlDp6UcScQBBUKSvCEN5D9nkxkwN2YEuMiSRur1sUuQKXU74jK6T4vcm
kbf9/tcnIqShMRYV4S+C/TPRxZmtHNrAjO64vJtM18JyDYpoa2+Vd0v0/G2IW3Sf
thqBJlRF2jhMOBvx94RUx/VepFwKazSLbzBtbzLXBfAEjVnBUEczBoy2zTw7EfMV
Vogr/FFU1nqix7GvT5s+mtQ6wSBH3T3V5UDKtw8ME443SkazmsejB38ak5wCYkK0
rJyqcwWX27AdAfbcTuX2TZnqh7gjkKh0/H4gBXARqD025Ivg/vaE0XX2de3R1Zjo
zlKxRy1NEdXqcshU56d4RJIfIz2oYLvzQxoKctz9SlPm1usz0sIVeIIfAWgJiP68
D6rHugPT93WR6WJ6a86WELAYN1y/mOhuVJrt7PE8GppJexoLrCsesU5NpEKOhxs/
clt/3YUUFo7R+1t3BZQh0ghVAo9qGmI+WQxlouF3MlLil3KBbu2QZX9swezkd4Ir
BGkAwNfJddZkN+wUY59QHMBh0BLNK1bj5O04x3+SeQxAx5JivsRM4xMKI+NWHpCQ
UW01j+yE09HK/p1NBDixYvAZyspRgL4X9bV0G4v/fPRCiog32R52DutsGK0bt4UC
tHbNp/mJgirq3C/d3hKOxg/d43Ti1yax59oDOxoV0E5C5kGXINRoUngzJNMjpFNq
ffYcTd0V5mvAWYW5CG769f7T0kRo8093vxMwC5+opMY5bjOYmhRczC6ZeLIZox1B
kuTfIa+OG4RZlBsUzMNQzDGdWNHskAb6hHc6n285tnxgY/7WXPdWESSDypYPV3hQ
4mmO0/NC0rgRh96e9omlwlCDRDUOlw203NXZASINTJDMaJA80Oq34aFK6QKTviIq
3FgluBHApm0PI6wmvd95JwhUqrCzeo5UexkLEn8ZTNH2if8HxWkkchag79HeGydf
fh9sD61XnRwBwQmL+hWCPvsUWcgXuDRifaeabwvRxL2Svgc9eIZkQh7vsGBNQGhU
ZWePOMB0q4TYuSeAT9reGOi50uf9XbeagxZOKutVMwmBBJsyGYsWZ3BzItkcj2m2
xUnJRWrOpnIJrqxwjN2UKtghJL1Xy7RtdhRm/BTFQkWx6U1jArosyqbScbq28Jy4
NjdlvaTXV5aD7KjOHWb21T/U2yCEhNna5hlJdr7FrVvSAMu3n6uoOCW0p5DNZzu3
weYo31ESKkUBE4eiXIAu10WR2CAn5ysQa+AS3nbtdcMnnxTKpXyU/9pAo0kF1wso
tGVkx723BiEpqgopFgFlZuwAWX71Xzm1WdCMSSQupgfuA8ljOtFFLPdlqwPbTQl7
S9cIUiNCFhtUvJtBUZkV17uOd+UIjoXQFmE38T3eR+iiw0bWJa7lcaaDvhruG3cM
aWXbVzzktoeZmo78HigxR38PgaMNb37JYE6FPA8KK8BIqZJJ9bGAFEq/ZDCe1zx0
7h6XtKhFiXCKbJ7ufyefruF80Q0RmM5zfS0CzUJGbesHvFDVjkaTWgY2wJ3HK4Yc
q/urXJVIdJSAw+fWx8uiakWA/cQHQPTJYMOxmFCGrCoHjcEh+j2aHw/l1PVTq+Ja
I9D8dMvWmQf3lBiGhJWc380ifK24xLwWqw5loPU9wh3uHxg6TU0PUVpNduIJHR5Y
lSGmidFA6dinOYPI8D9DX0hQ3v+OPncaP8Dtj8TjiAkYIgsAWo6Peeous8zsjOmJ
15e33LvZX7S+otT8dieQsrYQx+rOMCTS7OWJu47w5o4dcmSbDOwZITCKXSeWcH1x
E+RkhRvyd31YGs4T555oAEQNy4WQY3xz7c+/r7BZZKYToohDvnLgIqddNloTKLTd
/qrLaogJTx+82e0oDtU/5gc/XBVjhT9/q1A0+ICeGVYP07kk1A8Ag6U5U8n3sz7j
YGMWo+b/FL710/RSx/WbEkN7IuCJIz/5XbCbsFPtklQS/hABQtcCeAL4TeSknJ6k
wL7ED/mVUaCUlcoFm/4X+UmEpmpaZ37+IkEnOuyqep/yeoqKxueJBRZbc42GN9qs
WnZ163mL4sg7BxvAAJB8wariPWwdwD4QvIQoKGBGHWh5yr2WZj2uwYo+zLYjKLyk
xNPtkfbfjoo+S53gANdht6nlWaxh5riUewsGtgxbrksKA+4t3OuoS28bwXuef8CO
sSGYJ1CElwcuK5JIK10EpzK/Ye5JOxC8G6QOZsLe+V7V/p1Vd3Vx/JdyXPaDyS/o
W5EG+p6Vtupw4G1zng9GBcG3aKbTvoKxLOiNqJLgdN/sAkKBrA9nqeMg0Kdq9dTz
hBwTYgNEIuKCZ+5gsYeVYwWuZQdOyl9RFD5haR08L/QspXO3CKO5buBPQmtflpzI
FrD4MttkDDh63UtSm52/Kp8eVkmJUTp7pe3XgYRgQWO+yOpNunaOxeDx8KH0bE6V
3ylaK/h9JZyD3CtXgYpncAs4VmUUiisx1TMyKHdZTytsUKSKuBoJKaAiW51qu59/
ZV4qvsE4A+ZzyVWsCyE2QuF3k8dbsB0ASkrM9HxmasuZh4wd26kqoqpfqz32CndS
EhSwS3xuy5badDyPBmhzp+XWV2XRATSrHDBFGFyp9e/+VMzSEacUCeGuROsvOnLD
lfsycT2HwU3YKHeZkAC85SMfEadERBCiFwJlTPWO+lKycSzWePBXmBWkL5r1j03J
qph0CiT8Sma94RL6ODMv+q+dZmnXlWec8vMYpqhs/ZJ4r2+/1cIRYgEEb9kDZxgG
Y0v7ef/OqECjCQNosUWgmSr5ZigWcfkqu8tbimwYrO17qwoAp46nHOWdhqDmKl/S
E8ylDUriHB2XL0MN6KqTtFk5sMk7vCvRAAiJNWjDt1nRgKqprGUCPbxCJXDojcNf
QKFJRwk52FoceEAv8bsdScIDuJvGF2XCSjcIQIdo+Z/k/vdBZREa/zeoj0x6PCOE
Jw7NinjXhW2dyrjySygueThfZ3mAJv7eIjB/3RQ5x3ZFnFlCSbKnpBhiBDYLGMO3
EPEc7pGRIP4/eRocNfUMNio0jzws6xLAsREGBkybCg+aSv36JOvrDdo1m2WzSQn0
wrcwvc9CMMlhQIMZNKgbUQN6e8wWPiA+VpPwXv1vYLKMRuPzp1DjKVp9wVLCrF9u
/7DrE0K+ODEnvCycogHtoqVdQgWZz/YgLX/PC7Y8E1xtjbzKQQz1T+QT3GWJkLvu
zAMR3812xElb47W/jwUuMr8uWsUjg/3YgA8f3Uuzqi8=
`pragma protect end_protected
