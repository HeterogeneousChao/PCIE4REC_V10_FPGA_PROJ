// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:19 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L4xpuO1vuEJKtgl7AkBrN40lC5t4X2NKSnt0MzFHuL3nHZS+OrO0Vvi95ble5cfe
MM8R/d49V4xzNc1fuGOfYTCQLSBLjMNCIpjrEEEgx9Qk2qXAXjaAWBOmjF5dlyEo
v3yLuBG8extNNdYGf9UZ0/8YlfJ8wwcMUa0vAk1Gu8U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11328)
l0/3kYzTPX8XL7uZPt9IGSlctjuK1xJmN+SwHpQRnP749QBsHhqs0KZuzusDcnU0
mu13p7lIXUvX1ey/CGKLvOBRdfyQ3OCw2v/5L3DdhH1qvDrN5NPakJbfow2+TXcs
qtR5PIsqLcRSG2gmnaJBfP9HzEKNtgC5NuD2FQainKBcAaeDdoR44okkMQ/i+S6u
pJx0jDyeGDLKl7DkG1HWUdxk7sUGOxphEtR2M1S+aHdTQkVxwF5922PLss1u6Axk
2NOB3jW2FPd8a/5EE5BwJ39kRilXoJ141VuMZpCtXFt/LlWPRSxDRxbeLOYe/dI3
ay/mJc4cjR9zVxG2S22w4AN/pHhDwL763uVNH5wq1+ryqKD5hOLKJX4/bk4MJrN2
E+P6MamxnZIrIKkjnjcUcrxlqp3Pw2evu0B23LFtBz3BnYldmAe0ssv3CEo2v5ZB
2oINMDMbeiuzpS2oM7Sy0UqfVDMmLGpJM36b7A81VHXOXPojuh0URQGGz0o2P2o6
TUeN9BdkGx/+hQppMWz8lx4C+SR5zvbdsFjMVwvwYb0CGOAM6pxnG++bY0WZxNTF
cyC+L6idKS2aqR1OTBVEYq+B/u7Y0tLjk5N7hbQM+9+gv4pAylLLYJAOC87Ix83E
KVT3fkCTcSX65BBIIhp1j2zLntT6GyXIl8eU8/w1cgALjEei+rE7yK6g7c1VIBDm
zKUJXjbwKjxwhbw8ngLqUI9gVws8GUYfz/ckyX4Wys5nh8qVErM9j98+gPS91psZ
ANIys3P4YpN60+RrhmiIBV4Yto6pQeQKXInwPwB9LDJDAbPWE1qnGiD07NhH2pHO
q3vq8N4j1u61XcxhHdfi44gvmmcfcKu931MZJ8kXzPrkt/1Wr689zpfPaARU6+2q
4MWgA5VJhKkisNoNaMliZ5qoTwn1bTocd6TFuoQlvWQ+Ke3R7honDb/nMmN0tmDo
CWQBlDeY+OQO8ru0I/O0Na3+m+ePukuDAQ9Aykw29HbCQtAJ93PVYJU14ee90mOw
WdaaYACIzQEGKkgD49ZeMLIkzf+prwVA8DiiZkWCIejkkL7IB64hBtvg9sOH2Avy
LXABaW3NEq4NMxnEVyY0on177UI6sVM0e2E0dWkD2fJIs54axT+jvscoXZrCdmt4
sJY/jn6Yj8/++zKOLHzSnaszoTPWTCvnFXl7Ax8OgRcwi42Vf8JnpUFSDm+mHVJ3
yweclx3kt8S6gy+c3NJw9vVpT8gIy1FN8BUD9ADLaARdJT+fVsHankTnMu/R/DeK
K+gcqkIgxF0EwuqkL3D7Xz8QQUbGOS3hd7leYaYxnPW8hxv0iDZ7l5rmb0IYo8xv
DNWWN/3qr+stHH0oL00n9ehzoBiiRyKMkinWPRFrLFCez7Wi0WRALWC7X1QDm4tD
98AGU8V9igyrUBNv0Y/fuy6yMCE5VBFkPd9HYMayHWJ/l3sNIgPiNqtiGRjKajFj
4FScCtpmOXB9keQpS0Gk72JLRJXGo4lea5OqMIruMdW9+0hctNDGsHVytWkAswSB
A6mEtb9MORsm7x0U5Jp2Nb/ev+GQpyJUd0L9KiCS1orNaDFBg6UPDdCoMv/o/FlY
VsJCQNb5dZSmQIbD5MC/LbkhZf85s5zFktUfuUO0Xb2fhlLbWJSvkzkHjtAK1oJ3
tGpZp+d5bmceGZVrTCM72Wnjrqfq30ZIPuSbc+i9JvIR2R+Ow30nMdU53dISG6Vs
037DvXDGkfIh68jlbgymevgerpGNqex8HQ+lniuLBnLgg6Oa3f5MzjVJ2eUDAnhm
R3RWDHcI+YNbIShiT2/4aCdYVn7nRXJT/vfWtAx7DEfAdgUrXIGXCYo592aBtJCY
QXaWri4qe8tR71DIsQc9Njrq4KQAS76gBBID1dEw260ZSlOmYBhYpuCx9QZDKJGx
cALKKS+VU4gfLyxTXwKosSK29UziCEI2+fIknTVtrQmvB039/5MLb/tV/wgHXoDD
aWIBbJvizFplBRdtlDHQWM2lIbbSLLvTebafjkO+KkiplwU5ev8baJbprwoyuO8M
gpAaEcpcnN5bHh9KBiFto3LOHWCRRQKCNlObqz2Q+xxRfvIrLcyJQ4EM/pU8Cu1D
Awo23p97RgGvjkgGR/BCalTeR6vzK2MubHql/KKlhXNgqazP1ehsxgKi96dRMJr1
p3p1BTy96Onf15YwlvyFAR3Ke3Q/X6UjzOmbAk6wR0tMq5JSDELfyJb9J+fMDBv4
cmnQDEnX63bBHBYJOJot0XScgnVi4HrEHrXevVMeNxe0/9+1pTQT7Zmcys66cfpU
u1jajb6r/hjBAYOV3EFlkjfdaVUQs7dDD75O6bsE5+mvmYeXH7qbNyX7pgXpCREq
rWYsl/wpAN//jnj6N56hIjbRvFtmX+gpeTK6NvKMSa3e1jeHEcmchKEaJIIgNABR
6RgJ6iOyqoMpwt6dVoFwoBPHqdFPsOzpTFAGV/uvEXPWSsW47FSB1bh2J+TO6gjq
gMbbQDAh/OeYb1qYhNc99/xyisp+NRZa76BNhN+hiqs0K5yJzNlM7UNeUqN8DaiU
+4NaAd94rHOyj55HB4y/7aT3mzpVJTOSJxhVwkZZxyo2X43nqZcAImCvVxqB9glr
+HUx5PeTqAF3u4AoMrQspwE3RwX5RfuYAAeeogf0G9Ev1ZXmnfxjl9Y6Lax+2kz8
P2Ku4C7UzVMpgRYC7bY9XU+Qv6zIWnqQtKe3eByRQkOyikkkVi0RbNVzuLafacdw
1Y559TBIockGHCyOsmY13608RajyM0TO+c6vgWIoPGVmG930OOFNvBlXJtnfHCbH
GrMUnWraZkhNHAjWO+ppYv2o2dthDlMyOrhqL2sy7cTm8U4mv3sVA59ookU1xhCQ
sOmyv4r95HHozmSFPizETt65iZDdVp2JnF10Kv5Nj34goC6sz40aklm9GihCUSBf
k1GRQGFj/HIXiSa+BGcrbwKynb5yNlaYZeSPcEnpWFc9ay2CLQi8lIZshouPYbSu
tmAwg3Sv1VvOG6MUmPUglSGRrXAgANpSsKCp7UvD+zSp4t/8h3wZo0P3QsynrV7l
48ifpzCDQfRtFHRR+GAbsoCrTTH3zvgPtXbmw4t6QUMoqcduyTisbS5rNUrRo0Dy
YIAfJsfYFH1NVxux1pyalJAJo9t1zJmTpYi7/blc9KiSRIZzX5YNSIWu79cR+pfq
IH9UT/PWv4zT6wxhbo/ithdqPLhSPyLEE7+M3QnOzTpjjD+qNcONx+Hp+azUfWSR
LJWI1f17auEiDsp3dBF5Q/uJOz57zJQl17xS30cxuxnPFnEAe/pNQsxyYDp970Sc
gKw1zMYFj2Ucr0uAfWvvRhyU8tgk0Wxtlytr4jCLlZnwqF0XEolKXb3sCsGyEpsi
tRvYZcIZBiBqb0BpV+VYshhlOI2sZgiDnGLcIsSjrF00PanBdPtjIFbTxvj/Wx1t
dDQyz3tFqIWto64uM+0FZ+DVwYc3sma7IqBgH66Ahnmvo6CZK5Nmecz3o6pRTBhf
cgVV/B9USrn1gF2XgVzZTJtTfHngA50QhYhR8R6jRUQzw+EVXLoM8h1LNHL8heMa
YRHfXnUJ3pgfTwXWva8FL7iy+av9XkQitFICHxhMfO7KiYUka09y4Sh09frYh7ry
URSwHz5AEXu1jGWx3GN0X4Vr3GNycB4SEaR2Q6FSPgzU8wtbpED6S9xy0V4W7hbL
TqJ31B6cuKFZQkcBMXnUK8qJH8VjKFsQccrjnJaz1DN3rdB5QCjJwlqaJCbxWwTo
gEk1xvoVUFv1deMjOUJYotCe9nLICsZgUMVdRmhE8RHW4cFNOwK+K0IwTjILaJfi
FEdutmPnLVALBSPchmXJtowdkME0YHVz8evLo2QkI7794cUf9xYcn6R0e4Z92eon
8dqh6B8I32zj8WoHzGQJFUIXSSLwgNQOcls3FZTy8BX+1Af95Xxz9bKrWZISRixT
iaY7zmoOLAFyElc/Z2iJ7bKr78HNrwkLejq8ONGyYCjWmf6/+wA8CHtKTSWOJrbp
ioqwzJ89/m7swN7C7h10VzfE7Gycsy3uI1dxg4YmnBW0ziuVwG1MyNbgRtqtdkzB
gK5WTJi/y0PuK59CTdrfmX9y3atCAqSZaWxHxzqgnp9M4P2zJ5KjkUU4X7yQY0WP
9zU2JGdrxBOj0RCz0s7rHafJKxADZ92wRbte9rBV6I91lVG0EWOhHJBanN7ik6p+
MvQnz/rbJZol08oyGX1Us4i7gJ8ep9n+8SUmzelD709vEtmIXEi/3ATpSWufxkXb
AAH3Vcg8zR72OU55s6L9Jn8Dn0n6TJpEJ//05TvP84LzcEXYbWMgnPBrM83anuHP
x2xyRsQYiuFUx26AaJu75JETu6/Ksk9+wOCs/fTxd9ms+iYZYn0iE7VK5mgXLalm
Wm4VHXJrzCCt6MHpIRItxk0wY0wvEvSSRqsEZDCtVF91obWkDtCPt7dvBVQfuQhG
ofrBgmntjarlXR+kHUQhjTBbc8O6LKc0iPndpr0o1Hlwe5mVKsNncKQ34XO4jEM/
0cr6BOkI0gbwvIDJ+YCo7uda9SbwFhgMkFpL7PfHGcdatCD6L8y4+zctagMn78J0
rxCNjteMGoqJmmaBfQbHzgM71SUOHELfeXrpIuhzDb4cHDDAY0A7wrhqBLnFQ6zQ
bro9Twlab/N58X1JLFfOkLffenD+H2/ArVNPljjcMsdNlcSMJ2k2JPfrwbS6VH2x
WBDWOGE+HEsttWoR2kWZ662uGlQSLJGHtxvqw6nvUjtuBYvznuMQjItXIfOAdBkX
UiqH3m6lfMFVZFcHy7iX0FJAIXlJjOhvp32VeYN2FXjQwSK2uoyBm4rFUj6MWOE9
MTBcVDcPxBW1PdKZvPRqhQQjqrctt2nHbim+bBtptNFAscpGJb/S8sJ67XtFErBr
T/DJPijmS42XXloiNJhHfm4c/TdR4zdyYbNV+ByQEFmEdAnFr5AFes0jCOu4rGbH
bR43OCtM+D9sAqpYkPQNNIHoGY0sZdefDxvMA9hE/xPnIJDv/nqyWJmQt5mlu22h
myEGVgzoy6lug4/cP+0eAKDcWO2nPec+t/JlqAkRdA2ICuZ/sbp4X+mgll4UxkM1
72dzOxzABVDVEkMLwXlYWbTKn2YzkJ9ZYdKBa2fRqndSWsGKgU7hLi4o8xSKmKuf
mvkgWyIOxusLXqYEkJoZCvqlRKnCffcnW9ScZEEPmSAJpjrR/dhW15iiAkDY4QhR
eHmOfpuFl9Fv9WsjoA2jhpJ6JPdT1IJzAA+KpXZ5AhJ7d42xN+E5Fba4uCEmeFRE
ybGdJcMZjAiYKVVY+5cDDqrt6CiIL2SgWQrC4Yph0t/LUrFsR3Ddbidek9nmSjSc
K0QColiSiQhtbLrXPTYMXNKXCzRQBPJitg4FQEvXszl4rODqruopfQf1qNGbtDRm
tQ6FEJOOZk+6DjXi4JKLH8woyMQYusf69AcYjX3ISJocBH/wQeJdqJFZOPhx/g3k
zLFwDkMHoTjo7hPo4cTIk9fIL5LguNakNiL4W1HVanEtdcQlCcAt3iy9GT05kt1Y
njNV5qvq5v8ANhyzp/9gs2mkg1TzKzKq3r5QxIV8lPz9n/q2Sp9kydh09anxWL69
DX6NpBb4P8zSb+1KxvcXMv+LIz0MRrt+qWguNU1dC/pr2LL53Wb/jFIqFMLJn+Oq
JjlXHRMzRjIy4ux3uy6W6mDFMJet0thUPEBccrISLD2I2+4BVF/VMFPgXW7oZEpw
b/AXoUxdONS81qD4Q7z2Dmvax1uARz/pnr8JCHtVRQkCaA5uSCjyWVHDjTuhz8kD
J0zVXmjkda1GeTRwERrqmaWVY7pospCOf91INEi+tnZ8oweqsF3fWHt1xQSkx6/E
R1ZYxqYo7Xdugzg+Fpb1QfxEupRbtujXZRRD7roag4WV2NWtO+bKsAsMeJf//edR
gmmgcvyBCjdzrlY1Wm/C9aVHm69elQ9KyQI2VTyaSXlTOhaZ1kDBt0+JQYt4g/A9
38nMasdy6z/uxgbJcqmkkWLslyauJCitXAKedDl6mva4jdIUq5dA9xCeCkMqTQtK
KBd+xLfi7tZ+LlLU+3egehw/BhLQN8aoktkR9fZ7JUdhLQt5o4OyU+RUHMz9FBQX
HUhnhqI6m/9wFWVEBAf39nr/vusbM0hcp8784Ypsqibq/+TlZc5vuWeinw4R1hiD
HWOXAagjTnagiCcSppGvujtYy1gvoaWNrO744av+res+bNSXRA9jlPlvoLYPLXUE
nIAtFwmZQqD2YY6ITu1DX9Qn7dEbS/lpzhDXTpU/27RYTg+HezfKM2FpnrcbwT/g
T+C9H0dF+aGJ6UxVufxQfJucRa0AVmqUPghL6y3osS9hRwkDrJEclLec3LOjgP7Z
aEtwx6q6ESFr/UvCtw3/ywEjyAeaRXKBD9RoY01jDJ2fHqkNxXWRNyupQwuX1xbp
K3+ccm1hQVRpg2mGk+uS5tJR81UUWjoSw9CwtpPcg3YQ01X8jJzweTbBYkZnHkc1
02rXlN8FKJ0mB9vHAmVom1fu/4hbcBtrZ7PAjMTvF8+1Buvd5w50ypFwZqSMxqUX
Wt4kjBkoma3r01EzJ1pkMFuUls7RQ6GxNoMaOgyUu84TwlSmMdEu3tESgEdlxfL7
/oFwobayqHpzVYpLvyi0yOuB4GtBL4vup6ACOx09cXEp4930QgoyETFceu8a6fbL
I6u3OY7evj2H6c7HWtwJrWiXw0S5rCfHspcvksobTePsaWOprLxqZsJU6pXl1AkD
H3pPnKU/bY3Zh3fehlbsXEsxkqAJtM7+CaXfLc+PBSN0QPlYIAEgmPt/lk0EREPs
2CCO1QUkMgmowb7Z4suEyoRnzw0if6/XwFi3bJ/3VVv1Bd/OetbsEYd0HItA/x88
0n+4wlYFCG4Rvym0n1vzihaKMYNIgx3pOHbs69/za61EZFFPPKv83sV8kx/qYhZU
mDTnbAL9pJh23pnip3cNtS816gesB4esQ6nzMKAS53yKP7Ac6fZLHOQZEz0OlVmm
r6Y++xpYt4O1Nzi/4XEt1crrgppOg6Mr/Mdr/8AFsDFo09Zf5N92VkDGnK60YH9U
hnw1e3FUeIblRZ81rk5fN4tBh6k3rCLw8JZAyPSNZmyxMS06QAUu4yYbWv9xLPpy
jWz5wIt5yiihqAp4Q35tKEHRSbcOuGoYxcxpt3cHC4MxuUlFb5Bshv3DVAcjlwk+
mB3cQaThKbVdLilXYN1zjMOIeeT71oFZuqRSmMzruduXFqoza/J+GNXGQLoYCxbj
1SOvth+baY1ip7a77gWomsBRBhOzwct7mIehWeEKwykbVA2ahL7Dh/sYtepTEy4Z
XmWlAgPWmHjxfx5quxKdbQzRDMvLi+DaPRlfocoZxx2D6oK55zS8rGNtOrLHlSv9
Xi5WiVyhF/l/4m2rehkuMmtMLVe9mHgWmHJxneR1Bkv7jG5sU08+UqKEpoyfidBz
BuN18BrsnrCGl5QpFr2OnBlt+HJN8m/357GPuKuTi+LEtHE7zVEnSj0mUQw+Ff9B
qU9OTJkoMhY2nDcG55nsaJmzr+LJYNOAH3H1MD3tyLIyXigHDlOhyZi3CJlZp19W
RhQMsXqRc7zmb4Fe/+onNSw2CRPHGwFYuS8KZWdQFaGeCTR2xk1lbXXxySpfbKa4
+/d7A4CIzMrz+s0riGu2JI/sWPSVc8TiSmAvsfW25cpluHWSE4TS8Et/R+kO3dHW
bSZ0Mg2O3HOAbfJdgH9f5ZrfYiymooCULBixmNqO3d0FKlM45Px2DFC24yb7luFy
NpkIKLbfCfJy77RDr2MfSjIqv8d6xNb/tInzgCq/Hi6Y6y/6JEFsP3khJdmK0F+5
WQgKxGylcrCcM8Xn7DMK1ByJw1jcP00fQQz2pmXWqSUyWVNchqMBNXfvytZ/6cL0
Fpo74JQR9VEtwwMFu8reH38OSDlF2+VjiWAXQBtkg1e9iDqp8CtkvLTOtJmfDKD6
QglMSOIsM7ZQBfdOOpzPFd2TcjMa2A4+LN6s12RwDab0D97Ugty/bVbF4bl3teap
yQ5mKkRi+ozJ0u19V8APYoN/ENq9WxprcEu3iC8dHOLtNNdIrqstLUb4rXDXhZ91
MRQDIPaNb+6/H0hEvLKVHJzRzdmnMmyRs0l5dtWk6SVYpV+m932hDGn5qoiRyRXY
zE56BYPue1awZlC1hVGMG9zFUn3V3GZ8qr9HiZAMw07m8dcZYHa6XVQ9OldxtwcS
cQ2hOqb/wEduz05a5RW+1T4MiENFSrVAM5yOtUiVBXwC8Rhb3np11U63SdwqlOah
IQSmUzBrPHDsRy7oo2NcaA3LUWDfqJerGWupeke30qERRPSocb9KcuqN7SKBwUlB
u5cHuPVLjabV01kXaTX9y6fokGESth9KWeRSL/I9jpW51GM7gHDmnzp/L6UKvKls
1TmbtzYhQeBSKD5mEdjEzrA3hWVz0m6R4GwPsFJGfDO3JCW4Zo+6ajmuQ9FRYdiH
dCxY69Ew7YlbcSkOiuSPFt3Odjo7nb8HiuRs58sq81ZXj/udOLBybrlwWuRxXrLc
jcn8kVnvmOvtA9XDpR+kio1AXwZS0pQaQauP2A1Vi9EUSuTFJQa+rHYn1n2wGiag
Lz+3C84Mr4swO2m6WLazysEjt+A/eCDe3A8xQc21Q66vYo5NW9cgVuZH4AzBcoun
KQ7hNkR4Ql1f9R3k9afAwRU+Ue2hp/2YA7VkEQNr3BIHg6iZW1NUhhEOGsKR6YF0
G5deuUOl5DIZAVr835NTvnN7Y9N9ousO+tXT5a4UkyX+JbnrX00CD4XHndLZWszd
uNg9i0YTC/FgpbI01U9vTh0hr2ZC/SXt3i79P3XRGEiY7622UFfK6SJ44NWSxz6h
7OkEYH4Rk3I1thv4Kg0FTeh/f6RyLQACZ6ig7oRF+s7vxvf0qMwdBQnD9ZoEWE8P
3WA47lsntcwbSQgspWizAgeKoykfYBTCsZ4kuZLO1Te1nai6shQy+xAJGEC4HnT9
H9OHmInen8OWsdjXWIQIVDTigv3/VKdCu7x6Zcx5q8lJOeYyjaiTFcUdspH60trD
u/fwAPyC8mO+aT1FZWJEAvkZ064TlAwHD373xfxPHdNnS/z4vY/jU98i4BttL1bu
rlfOG9Fd3e9MOI+CmLUQIrs4Hie4wZkf8NPVZDUev1ruxbnCZVp91mvutnsoTvAr
Y/UpHFwJddZcMb5o9N5mHTPocO/d8ZpzeQnxHZxaSmoND/T4U+EksBJNCOW955+F
VJ5vB8VpOSfxuI8617TUNt/m7Jt0J88RgPrpTCcKvJVOONhe17R4UQ5MX93Rix1U
FW46u0O/AuTVObI5VvwZDdUZSILfhjUD57sfn8bH6ql4EhPNGXPIgla97MzLhYTe
2wy6gGgq8gTCP/6063HUpvWHF0g6/IG0E9tqSFG8TnVIEinXwrh3t3hz70309csW
9ng7g/ZtB2mJXZ42MylUj0yI5MFOMJMcGU/kq9EJfXBF9ufcOMH6aof53MRold2J
0ToJQAk5Wu7NP2GZM+NR4KawZlIUqnE2dVNU5Gx0jjazECLUPpUU8KuebWbwHTe7
xuC0T/3fVKlP1gyexTG9wPZNxErSrToiheDm7HluAePsTIKxFMVzKvG/+WFktRdp
WzygT5mfn169MYXbdkCEnIM1Vu/9TqUt+mIQobqzzInAJPM9MC+phSMmTSMbLduL
N4mkIEdvwlZrWyaB0ixUFLj2XnLMXWBBAYezN4jfBYma2+IJVN4fKLL6YqmSkaPs
fcWmqeWnnl/u0JGJO4wjjZjELjiEfy7Z74Hmq+0vuPg5jFALzdJjcc4FKkvwtru2
n7dmyohQNE3g4TUwnuT+4760dnuN/qtv+YqStr/JaRpWSrHAtFau8jvdOl4eLrfh
U58spR6kq4KC3to0stXwusXC7U1TdBX5KdUGBRJjLRCKWKaMZkvGGo/OgHcg1Nbb
l2GKs7WAC9/1TPGvBTBNepd5TrL4U9Setaa8El2q0Os8nwlhVspi89s4bNK4aP8k
acElly92bVr3tNawEl4cmgdPMTCMs95xzbVt4bqsS7qKfnXNO55uIHP3lS7guiRC
YrVToQdppmS7NsIOo4nIJ5Ljieu16oURiUOYBRHv65m+tblTsq4KsyD9/WQeBibG
v2U49A4WyC4Tx1f0b7heyKHnXiWDLjfSwb4nho3UKSROTWFuSRFIyYiTZhoFq/QH
2g0ERmjVFluL4B1rXh+vG1coM9PW7SOe8x6JZLfGzOrE2l7Hps/Ff58ZxAZNRqpG
eQ4l9j0EpT0lXTvUjjb3N8q4dgqdkqF0NsGTG3wMSFkl8d8PPEVD/frhs+CJvuGS
pHGpxNJwIN8YKMpyJLtFBEUosEbFL3rP5i2DfeRgyWd/Nk7W0ZvnT+UTwt3kdQl4
1N5PjCFgHZsDjuXHoy8Lc7h6PAMeD/E/cImXqBPyrAPMP3fKUmzZKjbPQ8cc0GHm
sfZtpxXTr0Ukh/6YbLuHpevVEDttq9WA+qwR39aY2jbeH3oPqR7gtiPWZbhUJYsv
oy8frptQFTsJYefN3Sctqp9Wo82X3N7aMwO4vlKhY4H9Z0YxzUn+MpnQD9odmRHe
5Mt0AiJ+SkJP/paUSpkzl0TF5RcNXCLLB05FxTXvZhVboIwysWxBCSO5oVPQXrRE
Vn2Nc1nnOcNR+vQQZzdhS13yfGggOnAzkjRHRAOBNfmn3cYZdKUt+Hw6T6Ii5nlK
xlSnhv0zJLzD8J+kS69HOhSBKP0hIT5Tl4IjupDP0V9jkgcvgFXMFanZe/lTHyQ8
KbQgG4Pe1LDJYQkjpVqVfcK1EZNY8JOYn8PuSS7r8MhTzt5BrsJetpvaLgiQRt2Y
IBlbRmh7ac18gyR5mzVsH46RYhN3Z4DQvTSmMNkZk8X0j7qEY76VJ3k/UK40ZlsR
NjIkU6nPuxGniuOaPmc5Q/+E51kqW08SynWxDIGcyu/nDuuu8KoyJmnXNnV3ajkI
fA8xE9iGNthoog0dJgvH1g1J3XL1xVl8Jy268+Q9GQ2kPAlODNn9tU78mQpTXFhs
8HDVBw6kqF0qI4af4uioUKVBdD5KtuxLLmNK9/ofoEEkRK5NE/jaJ3c0MMM2pKug
acXfyYf99EkMja4w0W48Whrb+7qCEBQNh8HpFx4hG72fadbLtqUEYaHKdowfu1y9
GZM9unKZAyr6/e7d5JDoIRBGlypdzWxFYrCr7AH+SBGrSiQbkaL8Z06U/h4bTaOC
0pcZ23shETUsST8niaLb/0xCT39k5BaXltLQ94OFD90+KtrQlFUaD/IwL55g9PaI
OwKObhb2CV9QLp5W5S01w+s9k0p0tiwBRjecktfdBtTBf9rhcNUvaS+rAL3wNHa2
8Q0m397vTQ4USiXkigfF5MwWWrb8cbsuhNdxUIImpjdBay4KrbAMIGCHSKTp6y+w
v6+KxuGW9v/n9G/odrmyKONJBNHOUpdrfCLYgrYyGslsWH5ErlSBUWwHeOOjCQUk
zvDJ/Walw9eHLIvbrJlZ7CIFL7VFQhI/g9Thp1SH0svop4HJ44+lBnJFVYcV8Bnm
mXxYSiQkeSZ10Ya14z0txBgR1N+kkPxfCLoAYctIFe683/KxlgBWWAAmUDK6sp5o
AEfixH5Mss4/4U1kS70WS8xoqmIBcZ3tI/EnLSQAf3xvH4kEIpVPwk6FzopWOeCa
9BloDA+XKAthovGvIOPYexDHYIS74RUYJpL5iTZU9sSQgR6B/MTD50E5zzXSjflQ
oewCJBFmuK4alGcc+JqI3RnyT9qAGUA0eu/9IRLWlVoCDvrzmrf0+qaxKQ64ugq+
+ndQf1K88s0qay35IpNoTivx6A4WanoBKehezOPaScE/2j+c49qxb5nBobrkKDfZ
g1kknrlVzx/aIGpdmJ48PRYnikHI7pHBkWEJ5xT3b/oI/hYZS0horS4Ne5OLojE2
A4CaiD3DmU2Riz6tqHpM3JWIUKNBlUnPzKCNZ+x4x/cU+JwoI7Cmgjtfzr30dGfu
cLVgoYJYoKkJOstA0Jkl4zjyP8UHEwLye3WNmGEjonjExpkt5zyfeGdO2vqMING0
TE5FscbuVX1VPxW4QC/KwVTvVQed7BrF86+zOvVYEh59KV4nGnxpfsUsW/Mi9nMB
gOMxvK30517BYoFawTaNia0A/eKDlQGCIYCJ8VskGaoCnesPhsxhd3lOfOI1pECP
KpZ+nvy9BKQLHHSz1iDx3RrBGd5GtGJ5htTZxDQpcddu/4xj7dsBYE1eVHZquKln
gRY2l+S3NGrAaQg1r1gcBlMG80VCJZ+QTD2p/YAWiIBebzBKD6/uzrQ79W3ax4tq
WOv5mp1PT3p6Kbu39fHW+tQvCv7Q3Ch3TF0gD90mriB6dgQH2HvVfkWtLYVaDCeF
+h6VBejH7QMwcpsiD9PHK/w9KhCAczEvu9Iy08apDbTtJfcjHaIDFc1wLPwixGZS
KfrlS/IFrGp/Xg6ZtJcOMQcvFDoILpoPncLJYzcj4S7bTnJFF0n/Ed2BILPOLsVL
lPpWstXX31G8ItY19uCf9mpoZvZbYhqk8EnmbNN8kFXsn5uHr5YoBcjMRQ2Gp5Kr
lp/2TW9ykGWnvQRjggbyvvYcWpesdTBb0Cq1Z+55QCCWbQCc7jWm+b9iOpoDBKYe
F3xcpPLtrm05reiMByvJ7F48Hn+zlwPwy4Xbd6HmTgxtH/LPORgsqvBrhUGvvUPs
1EdBYVQ9G0eCy4abybS9HUuPIzwka3AmPmXencHIZQIxhTN4cEg1QOxraLjNjtSc
cQIMcLBPp+nMd2fD/eS5mMNjN3D8Bej7XQ8nnv3kNPD0L2wMKjTAxVIBiSnwqAAm
OEtOuFi7z7/iJjv79RGch3DzRbOrdhiUJ6jvohBDiwxltYip74cqv6PR/uGY7+yX
zxNNVmQHu+hs5LHFfjSQ3/2H61PBFzVy7BppsjQRykCZPJw9PTfE8h9M5fjcEKCH
fV6DJ28Bw6Sn/XoLAhEZrgqws8DjeySt7gBZdDbamvwU18EBuaX6hhPYJlgMEO6l
kW1NnVrMbklliXLUZ/FCNR55JGPPk6iMGLviFF22kdYZFoq9cQZslPb5zpAoL7Oz
5FwrdnuY52GKhZJbxcmpBI4k1+QHXvvgy74hQRfDL+dIKz9zl/Sn2oelq3dxA0KV
SVzGQXUrzdzK9x8BaYzzjC/fu1BxFsSdImWzd5pZ4DrPrHmaMPvLDItxqU2UXFC0
NcGRV+R3IDbkHmJ1qErapqlx/A0JP/+VV25BrryHXISpb89b0KstfZhwruGwXno6
6PRDJX0+KLyZq1uY8/zeMQGlfapSAV9pqRFTmkT5bskYtqwQOaqwLk86zho57Lgt
mImSvYsPT3gz18cm/StTlECSTK/A4Nsq5/aT/iP2hrC+R4Z3TyxNZ3gUUkJyMJY8
ZRFFgMTFDAPVOgaTpju2g0To1V3mCphJLXbOMDfE8vkNQBsc/raF6G7m/R2KtSkn
JUAYCFiFLkuP5YfXnUrzX/tOzwbqF0bSgt6i3PD4qz1/4BTWonYcDdnx1vqyrGrB
E3DPu2Q71a7TibkPJi3on2DyUk4iLhdRIpCzRxBtOjvLxlL1uSRlOQa6PSuH4rhL
XLh7zvMAGHlY3WMrfDTQ+XBcs9nJSC7jILOftV3KLlT0+Fgrp/RAMOZXxME2nd8T
Fi9H8ePiyXsYi75MNXnZe4PbWxi5FkUYHPRfD3NrxXlf5LoDYCHoGATUH6l+wE9P
GiY9cc7mvpRFUvqTPshlhE08E4I71/lFMhaTw49wdwq+QY207xP4ypHVJ298kilP
0w9CQ24RSp2odD9livafZKwJgj/iUEccQgCO2iqbX9AxNOgDtFR1kudYspMvxDyL
WmexK9LE954dhim6svtpvCWWe7/aGQ4QrSnD+K6dwrUur/a6cLieUx86cLl4aHpm
1Favdg5BHqL9yOUBy7d+AeATHP1Uad43AvhKrq9OTsJWUeUO9Gwzha+5keNEwhz4
kXU0i2E64Sguik2Bbm/N4RBHWQCG+B5TpDghXmbSozGuoXkCMP4osEM6fCO88q36
/Bw+WFsmpSM9fpDiNhjblLBf/JVGaxqSn8tHaXzxbt5to/LlBKAvex7b+cmD7DwT
sWDEnlrAt6Xj5DqRQet9xg7yP82riBpMkjtTZM1JH3My0zhPILddGS69YR0H6FPy
+dTzs2lvS4uigGUwudlUQe6nOZozNoIP/S36eO3m/4mdjrli+WeJPfK9JXMmCnUV
jNWEGF7LxtkzVNf7XG+OVTk/Sy0f8FFms4qUi0w1dE4LNTG6URK0U2J+IJk8QqQf
UcPYmo5lVUIjpKX+bz5Vpzz9vPcDcED1RS+GOHWclqE4IJpK4S1biLMKBPOCVenf
p4pXTpUqjcWEYEX+jADd9jlyO7HfN7XtrPoCWHpVO06IcSbKViD6pu01HKh/Ir7P
dFJ4E7eTBMryJ931ZbLacfBHlwJi2M4h90Kw9ad0iUrxYlyp3s2h46yRiY+xTgMD
fWNaO47NcfFflM15/1bAqYhmopHDkFZ+6ICSUoCiX8b2RW5sM5Wnb2DZrHWE+8Tb
asnR+ZLCLuKDXisJ27Ogv3IXpbdld4m+FLFwT+n9TPC2F7mvBoQlXWiRwcmb0JiF
7ZVHFXwyUR2uHZ3hRa0SbgiE4Z8mRwmVulXnmANlMWSiC9CNxrbjJLohsQc68g9F
Iux750ETVt2QWVKrlVDhRBN4zoE8dVEAUOxQ1ruRgUZWQnCJxCDVhRfttVSlIFJG
H/CcsiDiy0UXX7e8jhdgXCsBDIiGFKeUMw8QqECQMOswd8GtgnoSFaSxEaP/sE4X
Ox+kjtD7M6POd8KHB2SQEo9sxI2AV/9xBkr77f4GZquN1XHK2iPh9q3SJjJMzWRL
U4Tvn1dhaplk4HSYV2FKr4a4oYEPN5OJ5TnsG10iKroIchMmszgVSCZw5srXfr56
RIim8scTSEdNkwnIlwkUw9xFeVIOq9dEqjmd8fLFsDRtA+769qbYh7qH2DXAX9l/
EogUkZl+Id5yNKiNBdV+NchfrLmBakTn7qnUNPKMpN9JdqI3qQKWG+1ZTausQ8nr
`pragma protect end_protected
