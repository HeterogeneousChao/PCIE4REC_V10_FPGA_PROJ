// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FvCSzObojqtqIrOIuJJ0Fbv0YAbuMwajZiESTqGPKECEWdRHoQiGmrbHI9E0JyP+
fPwrJLEcAD4SnDzL1kZDLHqf08JRFJUfwyocx49p6NhpKfY0sg2+pZlr6kvDscQs
OZ9t0Pjog7U1RUWEKEgaZrqTNzfsBsPtsw6IR9QHV4g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
vh4lX4hwWlCdP2vY4VDrwDOSVZhU6KrgAVfHlEW4I4KdpE7nE26wjBlQPsiNkqk1
k5Ngrw3VnGRjF/WrUiTq7zzt9c06mki3NX802dpX7nG6krdGQngYGdUoempNrf7w
kUw/QdmSM5OtB+mxXf+NR+HOkGv1w3La7TIzfDkG1fn6VIyCxGVu0m6oOdbMpKnH
SUOCCs42ZQAEx0BcJ2hqt3ReTO2ZzA/ZxOZczNPl5dfNG6cks9dCBJecGiBFAHx2
ZaiJegOu78NBahWgG8wPFI4N0n5B40VHWAM7OfpRrCufI5/2R+Y6XWBgVKKg3kCR
nPsDIY4aomUYVTmbgaD/YzeP6gxBFcrwh7rmIQ5JaxULflHWOVlRmDQP+scr+ko/
o0wMc4WUIa0oJ4adJFJkkX1kII3XKq+O7WW5Ifbl9FOUEnYQZnHUKqM0A3flnJ5r
+N6xkxpCwZsMLWmV0ylsz+Ce26dBG3g9v9OwWFFYKPyqbBr0F/JbdQFbH7MOSDtd
2Yj61UaOSmHr4npgeEd8vxvuxzAueISaz1775JujbpWPaMgOhMoDlevl3D9vhnzq
Q+HGFqKzFmEMAxYlTDtH7AZ9nF7f+K3+pVKNzKnOnXqtfujG8cT88IMH0VGscJyr
JhN9GTYgVItEknQObf7+Eq2XVM7Mhwk8xPW+HBvKM906aF+DvAm0CM5ZX7ftwXJz
F33c7H/Brw4fX6xoQc8Ez/8xXQBWzcl5EO3o6v/iz7O/qhI1QEFTmXVKhRe0A11o
TzLjNlzUQeU0yASWBu/3Xl3fwWtp6DOBNuaMz/TGykokb1P0gSmP7fOC8SfU6q2a
6EYpp0veB1Kp/ACUz/4+pFrxoGtk+upZAGjEISLM7Cvw84v+W5rnDR669J+BwTSO
pE0BYQWe7t+h154VisLQZbnrsKkbrKoThYWVPBWZdbvGsAFG/eEoaFQeNuRROhE4
5ooTREmHQqJEaEteUHT2z388BoaEsFCNiP4mFhkNjt5WtPOGoCq3JJ15I8LiOxu2
tay/wrl6kBAktrdVqOrfeMIxFCq8vOfJDP1HmtylNjTZfGC2lFzUVpxc/flgKZvo
0pNEguaxRTegDrWlJoi8m+KNrPcKQy5xmRsFNF8JFVPSiNfeyyLofppqV9TN5okv
ZGmFhiXoRQLcjscJF2HbNqAwVgrlweMnvbF++/fPv8wUEYZLNcPmXnZ1OkL/MAiZ
6nhQgruHmEe2bs2tsYdq0f7cHdtP4VrAJbEr0vexI8d77ZgAR2Z5QlBIaJztTRHb
P9KDdSqgRTroCT8FboL27Cmmes2oH10zA0R0E9PCMNn9Cf7+mmuttCuTQNe0N9Cn
j75nq2F+KPPTriPFT+Bgd02wDcAzUXvD7H9n4/ZsOt0OXi5PF8nlksgtjAzX4UYk
JeRhmcNrr6THyxyhke3+7nvgTL2QEg9qoTwE5r1YTfAJlNXsLf69MCTTpDB592eu
RCY7NEdOtjL3mOU3BU1AKoR1I9JX5EZiVixy4rJ/U7ob6jCXPkoS4JrhFIWxYybo
Gc6Ua89LKBOSJlrLTeKCI9vrIFLa6TYqVOlIqDVZHqP3sgKxGRGmA032rpoUhIeN
04Zc8Iv9qCBQ0JYN8g8ME15TaJTqL45reAUH2JVlD6fQDKWEkWM7vDBH5LEW4lCw
bw0dZzd09scf0IINg78+GzabzIC3DwTi10vz8az3GZ02RAwc5kftx+rjDGyvVI1R
JKYj0I/y0Qq6C25lkgKvkyH30TQe/SZYo1S7CsB/BE8xVWFeUnZGGUBSWX9+XyVv
JimvSUkO8luTOvAqyvRTol1lUI3zJXK6qFvx9YlFlpkJGYSYSFsz/qNj5fqxDEjk
/OXV1twaCe2pvCFMMTuOtn7VI7om+Lnzb2feDIbiTq7kqBWY8ojCbs+jxV8jIfL5
5Jm/lMFIGRNn6n5rToRqLEwb3ESQ1lzaVloa7GYz5PcNuUoaIf69FbINrNdMLL7P
A5Jz32TjEffcDtW40o/B6GeZ0gvtu5VPlMLpmWJdIj/Ultv8CCtbDHc5sJQn0zME
afWTmv9o4oarkjNSk21nQd/C4H1bmtJW51ciakCrx7j+S4X6FZL1kW1YK0pyF1Ms
UBOJIrlLz6S4gmycL7vKvBbIyPN88ft99Rbnr09ytSUvdULzokW+ZnnjO9+BrbcZ
cprVTwttWyuX0Wma/Vel5KRzxLcy1JWyjMyeRydNrWtLo7jQ9Hh/T9sGy018UC9s
hweWWup/jhOQ94OUT7DDNt857mU9mCXf5NWGPlUsnzt4dnXzRfbTpz6WgpoAG1V+
PqsNMwKZrd9m6N9lkX/sIBOgfKnljTtwYXK+VcLyyDbooqrkbnNgiL++wnKTpP5B
0g93x0IcA1A0rORv4L7veV+DFdmYzH42FwHNpIA1+TDIWBHsVYtu+Rm3Ef3nkIXt
L0ZItlFdWoWuGlaeHhuMw7Thp21GwJTpf9JdSbgW11nM+QxZkYSeo0GLCNyn1vnD
m/kIqmNQwCz3zF6vdca4PK9/BIqQN+izcnxH5lSJrXrjnWXNVSNXyFSDHIvFfo1y
6ODDXRiRG3xo+veBQFPwaea+KVhcZ1Yb2PgjZA0YVZjoH8LjqIFrAm6NRBWld/DW
K3gTaouq43T9WCEmpXxatHA03p5kB3SPGXvcvA+Lh035pOWku1atc/FHzaTSWacv
6wfzY8hf5tF4HjE75A1TYQNQPngzZa7JXX8MRNK9hkZWqo1tKf1HozEDWLDnu3/o
1EruUuTay7WPf8Js85gVORigg/cfOhg5BfRFSTIRayxDj2OEW11iXk7amHqwsPBy
o85aHJj+OmGa++z7P9IcT1EvBe68VtlqLHCBQ2NKb4ZDTK6qkOrxb/2csQBGCwFc
rszMC1NPBYH8Hz/e9TUyHkauMGkjfaD2KHDrOuCDc/utecJF+BTMuP7zQQF+qAaH
+fEYvzvTyZ2MrlqwLfj3FfT9Q6CImwz436St7V5rBSUEjue7VBujUf6ffYXfjRDn
/yIdTJ3eEggBK57BCLio2FrDTtEFGVDehDeMb4KYoafae80f6/Eb7gymNliMpr0O
oSglXBFzijW1k/YkpAuZ1Zdsoodl2qxdEJQaXFEp8MNjvFqXbMvt7V5mplZCJAK6
A6Eewpy8a6MS7oPefRpmfGBdSRfFV55fc2NfbYoB1IrkY/KNwHJRL17RSOgOb9uK
FyHtXlk8J57KC6AbKpMyBQQwKQQZUoE+MKcglXSCgo5WAMDp2kmVG5sR7AS4sJQY
kgDrZ2SpEWbloBcmvfvwlZO0yLkUKWxWaWUXAbNOflMZPGX8WNT6lO6PXgTGdn26
T6CKFpG7baHDKtxKEDmYrsSS0nfaLyD4apInf+iXcnqvh74vbYtCEmj4tvmCf9mB
i0QsRsSogs440bnajszbDB9wjQyYoQtHJuM/ZxWmj5c6wo77bnkmsWyXXhdOyERT
VG710Jxqb1NqO7PVOQFx04l0B9kk6nhgjQFMJXeI/sq4ZGadmtSyRaiUDTXSiRCL
eMO2Cn9zAOsYXv5ICVaNEPvl/9HyD63N93p45YWTAO8qbl+vn9oRV4B1GtfAk+my
2EebKmYqPFCSa1YBfCfDrX5kNjT4JCg4nZtK8i4VfbG6uoxYJHEUCbMtQX9Mve3k
irlPKi2aEaGR283E0fgHyFo3UoszoeyBtbG24//YBeac30ncC+0TsB9eTc5uevRq
9OVZOpiAFgpbJOn59rPwn1UFwl5MybSi/1t4pGH1zJ+2IJQ6oC0nsJ4A8XH4CP1O
2jL6D0hzmjH0F7rQSFk46mVEtGDc+Zxj/ouSOaWz6OeftgwWd2vmJlYllHfSpNg0
SxmgE/gedzEcFtCf0JiO37B3Wm5hAh3gMUJBOl4uhLy6SdtosUPCZflsB5JLjQcm
SgEGY7A55ERBbo+8uligx7u6QhjE8+ZsT1Q79O5JL4HR6VaQkuVkxmgXobDSizOE
Ht7+MJMoTFSlQHEdh3D/AtCk0zOHvYCcOijeA2bAPHrhTq4Tc3orPCSxDfh9gpqq
/W/N8fNLU8nuQXfSw6XU7rbtENqXqSzEvdt0tC35v0N7boGJfYhLYapx8IkaiEP6
gv76/r5wreVM5dbrDHKRGZSecgjikuXJCxZH4thMaCBfNOvsTAfH+JIlmfmjSB0f
qRy5TtIRAuvsLwNtU7Buxo4/PGp5Whjupe1e/NLdIC30ge2EOoNZce3EUFmQrgcS
uBXpE+SifKiaVYGFCpll0jJ71gUgEi0YlDd1nrF8hLfDCOVGITRUAeLWVujy9LvV
uPoh+ed0F8Alng/ADW1f394tLqFODBqqaFZl1Yy/Yn40uPfhZ4vATc49Kfn7A/t8
e59wBXYgoyRdEm0bxPE8EqcekmTHcNZGpsTm9PqhkB77gWoqRbOxQdBojPx/FDoX
LTnny2pbNbKX2kJMBbYd6wcv8Ew/M31j9hpefJ6sb4XbcR2pYScTYsJEvmx8nI48
bYFNFGi/aZQT7Y7qgExY3msNA3Wms8bG1F++OXU6SPwj16KIFv0oeTKR+Byreq3n
sgJjC7sdJQQDFQ6daagn5Cmh3AhyAETDwVF8HL5eqCCjlhZqivMgKclAsipuq6I0
hsknQTOBp886P3gQB524N1VhESQffV10rZSji5J+xYULeQkx85zWYi+pIDyBTb2e
fBaEOuCUBVWXoCVvdpYshesOIMkD5pcFIzmzAbyFqyQ60zRaZoiI4GBpFFOx5VOY
ZP3yvmGZQ8ne1E58d0VmuqoVob+381ZPuH6Ri7A+XdREmEyGtyUei5S8EZAkSUKi
SSpIKrpqu2MTzpARf8xik2WjBvj7HGXpIG9UTI4Pn7IOWw6wLGeQmJuTutMrec3g
5dyI1LUP50VKWV2eSmcdIvDEMxW4swBB/BNNHAtycARr36On6XJxFTvfomptIuQt
c9QYbXb7slwmgYbVuY6SqStbGbl1RYiDZ2f1HsGAl/R+YFoP3ZzRX0SegpLhbdON
Z3UjuRyN2Ngu0xDzn4rUi+9X6P4n6/s023zqU34iIFHnY+DunJnMA9iiDQ/sItMX
sPfovWTl2NYudf8Q3J75y5mmqB03uEpTke859nMrN2BK7JXLKLptD0JxEie+beHK
9eSpghtzsPPlPf5hZw6infDNvXBOA36TaQFxARlJ8E09Rf6ijEDa/S0+MCIz5v4L
aM9eVcNw9VorMWA7gO+kRTjM4aiqSSJU1rsSrMxLctAfFw2jFncUuKTela9NW8yC
Xz0VfdT2lBV4kpx7AQsKhjKdGksVkFp1n0rFC3iW2HlZeHQ8VQfrpLsW4J1OmA5N
ko2PcooWKhRMRy30kds6/eh/5/Ge+zlbwk5+II4r/bTbTOwW5ht5ln2v7Wo0tLhv
+nGlL31+7uEjXGqgLzrJtISzU5Rtn4IezJx8HjRDO0yyq0A04bVdUuHXkpljbUz+
IS85UuWTzHwxhnnwAH9gnc9cia/wi+njPPAdBKY3duS35itCd/lMJ4JyJyjW4mud
L18dcVUVO4A1D3MYAmMzlf0kezVQ+e5XVurKn615sPzyf0cRcxGQQ85XG2yfHhLd
do+Ig7MWS0SynadcLRT8NUrlw1ka0Hj7/rcsk0ErMQvktWsCqxpBLllVV6hSzyDV
PEM5ivGzDDKVjHNWbXlzrYfQxQcAErharyDAQ21QwWNFuF16eJaXQKUafHCXOoC/
kkh2W0rUW4VSU24jwinpumf9WlslMXv4aCvfzZESjUpAIeWmO1OfmKYmHQVIDPyM
bZuqfPi27vN2b0/qcnUCExErWBDN7kMQ/BVvq8h2aegR6D+s2k04u+eXac0/boBf
DPlBH4DvIl8Wl99vTfA9ziCNPFvVmgPn536752xrodNi0cnosy+Xcc6APcQER+vG
8FD1FZBgaK6FNXMKSSYXa14tnll/T967iNkXQBM3sA8tcCs7fxzFC6oNfyUKvr63
qgD6J1w6ExkSFX0C6jxfXyuqx1ZO9fGFEHGcXXYUMmPfjGymX5gReqoF+4fWuD9+
Y6TqdKwp3AYMHRCudSQUsVihXmSUoE278uuoXJaI9iTsiQ1YKWSwCW0CgvHOsMzn
CoS/8IxEWvy/FEAO4yHrRJ3sOferyMU9xwAtvG0sqGovnOVVnGP3AchCm+3XyFtb
bQz+6K8lytHeZ+V99Tcio45Yke8f2R4QfCum4V3DOHZWYZlRmGHc/I5Zlzt8WKi9
F7hi2szyO3AmRA+EFPEspVdN20KqelZyTJg6xDE0PraBfjVPbByMfuOV4dy7Csm+
9/QmTC8RHhBO3I571BOUuvN7/wrh7MBGyy6TnNGPnlkO5qgSgAyGq5OBVr1a1/ru
I/bv35Nl+KcvK93gr8Yn3Cp+qO0zvYUuto0DhtYrdQk+UWwWo+XZJBHtEnepG2J5
oR7BeRRpFbsxGSXkvbHgrCvPwtGwWqudZulxkZ11F7jjUAagiCdK2yDZuuY/Kxg8
A0DaSgoGEyRkGBQjSoTJiVaVsS4HqAD1eLOBTQlneySel+o8CvnpVX/ZGHuexet4
ddRnAGNx5esqjnr4wWHV2CvCYp7zNzi0UgzbUEE9ZfN3+G6pj48EsIwT/1NIpZXh
BiX77QMHYUU01hP8y1vyVEWq0mB59bvqpwI2nujPkY8r4c/M/FoneAojvJkeUhix
RVymYp7zFITB+iQ4iRU66deV78EWJcGhjfaySb87oApNiS+pMa3Do8LljgC/gOPG
ZwCXnRsyDiC6ayUspqtedzz2mgUcw2o3lnrUXWqt2rIirimHayO3G52zdAtqQuaP
9bIgD4xYicPX0YoCyF/ULFNhyv+gKTzWuHzDyyzDVecZYPHmBEYKU4kXCi+q8h5Q
dfbCfyVZYhYfxNSndnVFgwDUk6H8pCWXjz6Pj7kllW0OjrFU8mQ+sV/KDAMnT/NP
rJWZypanZjR+EnZouelIAnN0IgzHx5pgsHNbjYXJnQ+/ZZKa9Qkpzb3FmwbjBUDq
YZA4dk+3/TbRNQmlBzOabrkA5rdOdlqY6m0ibdeFj2uuc9JsyDC/Jm1tQFfeymiw
UWue+ahpXMMcOlauDqE91Wy1NCZu5rZ1A0R2PO4AfizOmCy9jVYQP8NRGrxOP3pA
g4QiF1CGRW/fxeIpD3AHPubtX3idpJKEtDjb/r7LmUYWanlh6i4b91QNM3HM98jA
2aOGVCZGe9SqhfAktKDVjUfIo+N1NP8oHp03GOyZw4xCeHpVKxIZ6svycsTL03pz
UDot4nrzNSeIh9PWIMxu7IDG/plcE7RUSbY9gxzKyouN6UDz2AHDIpxXtSK0teYx
mExgqUWceyNKwIoAorTPoT4hI9kZ6CGcGBZtpEZeptL4Fyo9EncX2mLb9wOwIx1C
hWJEiRv7vQlD6J89VWcG/PxEW+Trw+rgUbtCJPPKfLzdQyCHtsbhhwNY86vhfryN
qG3TuBE7tI/VqO8bTS06F9LNK+WfKU+fhWqJCC8OZyMI+JaJ70ZZyOhv/k7cstRc
6Nx2XXrlT9uR/uJKnikyeH5JAVdWGqu6cL2d9S4mTDSeMqWtVfv+59tGP2t8xmU4
g3nB83fRTMxGUY+dxmKl1cclP10Uz8Vf3u9LHw0kYe02pVoxhz41wu6BUNEGRbW3
WxWd6EHvqh9/u6tOoCO8v69rwxaUHtrZJfsmsJwW/LmeyuehFXY41tDit2JZhmLf
Orv/GdQ40Q6ABfO4UjCEn/h4S3HGknqWmWfRYDOFjbjfCF2fjOIDCYK9lspLOSLG
4k9B1s5uK2ZNszVNQzf+IMoq8o5SfGCVFbsnoPfhLDYhgx5SoIogS7ROkFMUioB3
bPcwyGomj0tbKTkPnPVQcuAyqTHAwyBQELeNLfvUs1225jEwzA3z5fcU6o7mwxVx
u/RNyaOVu6CPgrBhTeDSEjJCXUufBosxXYtA5/DLlXd9WeOkuUhBxwL8TdtQPsXN
+FLCbJ7G9+DdH36td2ae8R5ZCYdgSQaMJz0919wJ1jIiScB8SJr7rUMoKghBF6yX
yPDY9yfRpCeFnqvDYFx4FUuQH1QJZZlsQMJsZ4EE9Vw9UHtVD+Xf1NQ4zNGf2GfZ
VBEB+IqKpZXKtkUADfzFa4NtqFpdgj4NncYfpysBuepHn6Luc/qNnvX00/BsfmQK
7vofgcZsOwrcYRvcpl/1AKcrmo1BAv38xZbyRJD8/U14AvZFls0UFVfqeqQB5A5J
0iNnyO/GBqQs4C1lN+N3Vhd3Ry8kBgVNb7bC8WN23ma4sfN/zV58jL1nKJoYaIi/
0Ng7Txc8K3yh/29DdYzOGJpRMmlfsrB0g4eelorgAuD3NGeRa8a4aig3Q61hVjQ7
N+YgGfdKWB9XX9XcPH6Xt2ai99RjwYZqaG6QR77yNlYgidUHvpngfDiTobKfULDS
1C+TM1WM7AwNWptwwvAxkPnGlW+LnGrrHkOuiqRiYsQ61wJWJzgDDEAxpD7yqoe+
68vtay8OyoStr9E8YvH+m1t04yfq6K2Lvma/fibPcHkwf+o28CbKgWulCKBSnXZu
im2RsczZO8Jkp00zEKfSSgMttrurhi3L14TfNPJVnLpM5bM8yyfVWXL3KX5jkSdi
kpf9SxmK2KvQeVlYE7dQLAO0a0Q5QG/RakRVZUDyPqMtMME9TzvAgOZZF4KYj+fQ
7NFnFO97RQV4jEpNFysae5UJiQ9/FDm0RXbX+d5mKCaAabhPfjxdNtE7WWSUElNM
B8TDZK0OzisrgSI0D32Y2dUrO1XSWPVcn8+1txRAroZPXkkbhDEnxlKKbZ/XTV/y
ro4ubNr5u2uSUIU+QiL8m717oLrv5vi/HS5G2aILyiVrXKh/s0FG5LhVXP7EcoN9
vBfVe1VFvUjOm8VUCnhud0F29R16JpjKQ+3vih75rf4hKlZFNKnJl5aJqAOMDmhB
7Pk9C2fQ2ffbUOjikLATYUy1utj6dKpaYrkGxVz40D3RpANoMFXzA4AE76vYm6yl
hKAEmLoyR9ZoXSHl7s8KGRYAEmFwJguZ9V5i9J9xhT6x9WPBCZoIs8Cce8fwdKuX
JRbdwhGnC12X9BkS+mfkNdY17CdWmmSF1UMJ0mOPUt+z73VxsOSbWiy2EsSFpWlO
HEv/VCbz7/JxFPEbT+MHOIJmKCNwJjGtFaO2KPu5IjePfCRCf0IQj/CYzAoBI9LM
xSVk9EYJGXb9h9fMQ+/bhAiOq2s3dl62on7lXZvT9zw8arDODkSKrxkpFazBWMr7
cv42ztAWdfroiKy5G+U6kkjbLvDq98BOeprJi7csjw4gnbhwavw5XEWw+gb5HY+z
9rltYwKLyeVBWtkjeOY6EoW7yIEd062X54dVnI0GWD9lKFya5qIxoLjhqRz/E1hq
n5GYZAk1yH2QMvIINg8e20h7DgXW5487sIfIxKSQNnVe5INSZ70DrpHjOeX7I3JL
izuei/VahOX1xLnGHUPPvSYxrkuQFxWQMP5eBF+OX8mwiq4McFfDMpo2m1BQZTzf
XnY9FGQcH00QGTssNxSyddKPPl6gCq/YCXiW7NNZtQ9r7g1dTEJXCa0gPFbw810M
7x7t4uxhZs6LWAF9sXatQLgiGqCEdTodWSxDcfJ7WQbOK4jIzUXelqzIKJp2VZGP
Jkd04YQ0/aO01A3u4rdeKw9IoCU0pVSgFrdZmE/T3laJJgwx2PqM5yE0Z5ufLtg5
4joYRYxYh+LJiP5bmINtYZljZhrOc7adHmEA1dBYTpAr80uQ8xG0FWuXpWwgGUjW
UZBkPxIyhzxBqNd6fSA4zPtnV0Fe8NWgnFbzbrbdjZQlwLi/p1EFWJntI6EwuNCj
AmmYyj8mFUSDH6wgIvN+QlUlQnJ2wNy3SFd4GPXbdjvV4pqV13mDXtBL3xUhdC3/
+ANFn3BsQyQDi1qJbqDDylgGr3vMFnLMS0kG6UvHN5gcb65ZCcR2P/eQxFL16AMD
gBDtX7ZiV4/A/NBcb7psy/fEEpJ6l0Vv1DcehqolFOD/oUWyTZIpO16OkynTLkMd
yO/s/PtOYvVz9byggd4H4z4pAKyLEdZhvm54znzEC9BWEU56PFmBldwu3TKNgH7s
ILZmxELZ3D4U5TrK+TBM02HFYEG/7AT6K87ZTXz4XQw=
`pragma protect end_protected
