// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:28 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P8wdUqb1l9wRN8VYvVk4mn0jXUv1/131Ny0OoK1nsB8CQV5mjbBzGXTPK4hDGxpj
QI75zJfoRlW9K3UzC2gp8H+skKCcqp9M9zbSGI1DGq8WPh+LFGKYtASrGFPnb5N8
oF7L0gC7swOkYwysmip/FUb6nXecDbW9zNCWDHQmQlE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
gfwgMahj38Xlq4gnHK6Tk2Ak00GNAHbHdnEftAe3mmqaTi4KZgwRiF7VXSFX4r+v
ePmJusdLtRKp/LeNaL/3j/UBtkZgWO+6Jc+DiIOn+f25KozpXKqhbDAAxex8Oc8V
ZkLAnT3GFhsMj/qxhtmex+m39ytcBePZcRE7kAwR+j//7updiT9WQHm1RpgQx30r
zwhYZ99p/W/ajFOFnMMguBv2rIQAJHU4kT34cNxu78xrufMDANp5DK4itfnM2ZXG
rEG4QlOOH1yiwoQhnxI1vH1wC+KRq3uCL7zMW3HVHf8ZCrCZG/TXSvTz3uk0t7BS
fXwVR5mqbNgbTEIM/DJZQvwXLrGCLSIbY3aLNEM9nNOifijTb+ok2UhAHtmp9tUj
LePHbHdelFYCSaZx5kq0lSoRdfWSL86JqLFCag+mL97vkKF9XJpLnlTUmAQNNM/b
ECVvcpR+wnfzqu8oEEhMHqaENlA0wIVDKKkS1bJQqGPerQwaavu8YAQYS+W1RAzZ
zhZqnnDimM2WHnsG411MFSge0rIWd1DfxEHRO2wMEpw2UQ4bfikBhiqlTDNCJctT
js046WEEPR3GEVZz3HzQJgylHLut5+8XflRubzRv+V8KVWr+ld32rqrg00g/EUZA
47LBaC7hZs4XXwNvoRXCzXygwZ6pKdSSYbcpTquZuP5Zsc3D4UIxxDeCldXKVT0G
KUdBEw/OuImOUB3zmW/CjTYzcxNIBZG2DuAOpOMQN9ZFVFqBUysikL5UUjGQVA1q
8m7vHSaeLTzaxMWYqEDNgIcesVyV1PFA7WpEZDhScxLdiEEtzZlIPCpEN+/1EbGk
ozbsV9C2bxfBWOhGJc+Kopxp8kA64KBRI/fa978EveLbTtpFpV2NekUejAn4rx/Q
1qggr8dVPGVUAWGD7lPpIjdE8yg1xODQ0XRuK3rbyBTHc6/TvTjm4oWGK+N1q+XW
OX+DKMh4bP4FHRxYuqYyU8c0YldwELGSZrTFhXQcrw8bF4parz+R6x6TyGhyz1H4
0heydDoWDwoKmXq4pQRxWheic/V3ilTFShJTQF47Sa7eEfLWDLNPT/Zabe+Qc3Qx
Q4kp5NofvDxDO01X/IOzD+0MsZMZf4EEycvLrPqyZ0RQBFP4FWfgRIL7wK0hVHpd
t1ANL21au4L67LuuNQH/20x6WfptxPHYeHFQAAl6EOwV1vrNUaRsZaBAQuZjzWmd
wCU8OCuOje+aCcak21djxA4mYHu/wp/oipao109HpKMfsQFAXC9J1RB21CHiKAxR
wZmUn+0q2fqiTEY0bCKCNRosTSAURoti5zAP4XtfKcGI1mc0IX/r1OpnA/XZ5ZfY
sT2Aqv2Jd3/jHOP35fuRbRTiLAG7GjSE4nClGRihOJ+LRtO4qFPQCKdahxlAyX5l
9ieEQxgnFNxdUOaDcWGJtd5y+TmlbhbAKZDP47zPDmupNJSX9WGEna6grxHYXL7h
QqQl8u1rMZ8DQzqvw9no4rd6hnOYDTexzCLlxyBgF0kgnToNcFbb8oNoytZZmBC3
TSRAvBFMBQ1lDJREaf81c8a0aH1hcYHHRQU8eb1V2nbTxgHr8DA+M7Rrx/O6H8bT
0ProqBbPm+kI0L0M+hQo/Z0yxWs3mC/815RqKLnb08UYs8C++LvTVP2qOwNycDoV
2ntEjUcpPvdbGWO8ww2wl+X6EVE+kSFYQYKmBU1gFzBZjBdyWAICUFTyUWso7DIE
t9rY195JKvXtbR1rNhdum3Ro0OACzs95vYy2Y03fdIHlhX7zSL08MhUvnSEwtaTy
040td3beWQ7ADXVdiQEIRrXQDoTj45XQEgna5zmxesXhQ4hpfsbmSFofgnKvilZ0
JfvRNWOLROwx5qEv0ZSksp1xjWE8PXUoZznDFMOl/YaDNae6eXGQPqKJy/DfPe9k
pxikNPVccrFAUT3896t2q1wJLH62z/cZ77ReBGc9lxySIRPadnmN/K96mGEJCB9f
gpjOk2qzXuD/HEsD5hJwaKjLrvtwuNqlww/aOUMnwQtrKupQLs8imbLNupR0uEkO
VOhhi2PnsW+MHWR4E/HK0uaFMVihPQwnABLAmFQXa5OBrpw+QDW8yXOkaPwyr7oq
S0Mp41cv8akRa9EKKxGzvU3Bp4vsZozzZNKZC+/gDqWY58+azYOF/unIX1WLbgiF
ar7qRWObSatjSSTtEV9rqjVambr3zM8sTF19cnZNkMYGAzBLMoCWFBf7qZQ4jMUN
wkMbJ+ZJvGVW9Bj80EnkH4s/IMuqLbB4KMvDV9FS2Jph/39Uwglq6yPBBh+byyf4
mXpStlkdTk/uPC884nrfkboqYcW7B602uRqfdiiC4vtjvbkIu3y38XCrDzV/uwqv
OeEOerA/wMcnUME4no6O+RD3qoFDxyX4tOgJyCw4cbMKAv8BrwX9qSPjyxATzxwk
GBApla/HrcvxF+S8zHsVYrrW03ExQGCRyYQ9UbXr9xhD7ClcRQVmvnQ93NFzFuNP
UL1PH8i7yc00R0/gMNM93XAHlVvbkvfYAsMExucEZ3B8jQJVmYBGPBt5kVoN9YcX
1isNqgfk67jU7NJ0bYW85Nd3Fa7qRtF2CmG3exzzSkiled0mlhedRY3MLXZNWK/a
iyjwLXtHlrbTwaUUiMfUonkKR4XN1MACgha2UtzPkP6mJeDU2kHuPXLrNuVO3uDs
mHYfScnvZClEdFHpSWMtfTFVgVB24Fh+8x6Nz8wO2wUGCrehSk/bdaM55tPh2XM/
CgLZvYqmorbG29BCav+tvRXPP86zNsIzEnKebRqJvT3KjVanNKb0KiM46+/fcIqA
e2NfjIwqTSwfThc+Y09qPIdr9Mmx6LXgh1j70Q5ETHr9ogN4UfSF4XUszdWkq/mW
O4MI0aRCkKSbR7Zgaw+D/TtTAuN9jKIf7Z80Qpn8LJv4X3chJhvBYPtjrJfO6Iuk
958uLEFxV//OGAwdys+steS3oKDn32atNTfT7tyP44QnTOgor3xDlLssEMaq/a2B
vVpJe2WhC3J7DTh4DQv2p7biS3NZGAjukA+eIYb00bMeDK4QpxUtVSNwCU29KlO2
4cSzB+Efw/bqQda+U3agpHgko7iqPNpetXorpIjxh8dBNKXjdHbxgXSe7zShGODk
K+BvKcp+yClUzAmrk0vpxchrn9OjlvXEZFeipqRJVsqNLpezlTnDymYrHQC9k7y6
9t3nnBzRZDs69USt2pfpD4SZ8PEqhsrVwix4/Cf270jNKhtrvwcRi8n8hGWeQ3/d
ohTLaZrfEqy9sWqUmVf1hRLZ1CMH19j9uQn9p7bxk4bSh2dlYTn5PfGGWlxdsvgH
X4+uXKVlcVPg2hSQzVCe6G9LlJ6aaxW8YWRK0KN41X25LjHPvDZOqW+jdRSJccAl
fPvhl+TQn4LuduRtdoXpEIsuC+1yjRFmNecXpMPbH0WVp0bqNevGnb9VBZVcNdcc
nnpj4yB8esktLDgL57rS9k4qtlcA2n0xCdsbwNv89nmA4wOiis1NJ60chVcNHhg7
qQiejSdXCIHvSCSdb9PISZO4WEcRWSS6oRoCCPoQyWXYQC6wyZyrNxamD/ANd8n4
Ou/IuOjqFAySZblAZ7lB1+GLdc/ZdfKoMjtcy+BvCjbTfALI6GC2fLvu/fNBgfV+
1HglZ1M7fFGwq/EEuTN/Yx/5WVbgTeqNch8rEcqoYYEe/UNiMZ7u87gTw3vaLh9M
/ezjlkVgftdsxr4dtyQVBMyofns4bWcldXjBBzla8f0kZ3FoIB2Uo8FjHnw2SRKC
jp5IiTdbIKE0rVjKFVsJqbrrvWu4MR0Zov/DttOf+yZ25kJvbIs9yJhkDO0x8LJU
qWp6MWWCaJM4A8qpA41RcPI4zonpHbBoGF9hyHlAmgD+KAvFE1/m88aDGgFuIsbI
F0zdQN5boyMy/cMI4gS9HI2xXYUKGCkXGyOzOzJm5tqitzakyr35Puh4vVGbduVL
pEwlXapl0V9kN7HQtz0bUiu6fWUWBcMpdaspz1zh+O54oyZc2D69E2hpH9cwvo5E
mUkoVO6xEu49FQypjNZw7BfJ3VZ9McCbG7ENaoarmYBTA+rH2DogWhkr4llFkCXr
cXoZiDuD+GMWVuTME251j173GqHAlqOBrC4MsdnKBwK2MTYnlxl6kjyKsrHk9Bdx
1E+81GncGrqZEDKy2GCHW7MTr8E/cmHrQyBAB13f41soyAJ42fqHh7Sj+1J1IRRT
FnzBG8Be9Q9P76wKOhJzUE7OmqSrcVq+Ye3+fy/CtiwBxfvZupLEbQOIAj0G3OdL
4J+jN2G3r7Q7LeeB++hHMp0k+zfF14+vTAxdBHxdRO2X+YS0woauIwGbTcKfLbo9
heVmbw2aWhhoNI1IK/znJEBmk18nFxof+VrGUmLPWT6X99OKzA21ie+ZlH4QC1tv
U8NE6Yki/H2CQsDZ9fhPynBUZOs9LAGMvIA3N15F3OMODV0I1ZuNtKlHuzLEu71Y
GkLIrICv3UquS0ELmr1q2t8VDOR3VYOdBO0iJhp4spS9bFljViBBP82WDdihc1uS
WkZfszB7+omWW6/mYbY8USpo4USBpRg9NB4mzXcG71fTlF3P2f1x2HJrhlfBWdH4
QeUiOt2clDKM+0U0Rzp6DsPyLDZ+fqUqc9kPSZ8GmG8EdXJQXg52gkAOUL3/bHG6
9F7/HPm5bVGVBHh55solXQBlTDEHJN8WF/jKvF/8S+RZ6PSxaMbfYChXzJv6awex
sKd/JQw5hHghncbeCfdBk+XJ0sIsLf/msGMPhCb+Ngd4TMbrhZuE+6Nes4CnMpxx
THA2ieLPBNL0Pdi7SOeKGcDd2jRWExWIecwbUqMmz9e4gwkJfkx467w9PGwJg6bk
+BVoW5sjZKsQvaxEqVVqMo0QO1ce/2r9kG4jIU4G0dM+w4Bw6yEXr1Cj7fum1T/B
L2Up5rcOZ9axvvO0K+N6SIKqufsN9BHXHoRVneNW8h+dghSsXNLXd0WZmCHHHCLC
7R8Vdkq1ZLlqS2iiGRY5+CXM69rqJWkJQgdW9Tf0SLv4CMqwbCq38BQTKnXUxz31
ZBj13LxG5igGOTQOtgWxrJMdrCyEpdig2nNcPZKeEg1HswaI8MfvlMKuFqRkcy5b
ATnnE70zQsmaWIB5ZrSJUutL6ij+I4rDJDpwI2ws3QlGqZ/R6sfpA5A+dTiV9HQ8
9R3EUB02k+yByAtDs6E0Xi/v6nev1SoWxDDLWQflPXZXkFyGzpXhh3EGQK3MsUD7
OJZ1ra2hdfqUVh5qdWhjN1oqWDSdETm1MnbnseeQGZ4j7wm12kNvX2N1FKVG6U3v
xGHg7VNFHQBd9wxiHBY18J8PykS1mMLADEawCjB4oOJuOzHJeGk8gO7o473R8pNj
jZyEXo4qZfB+OuKZ5FEGpX0xywBY9Gw9hjrJ08/KaJHARgd9ohAbcXxitocI38tb
VCZsOFnEBEo3lMK8DS1lHk6rWYs9qUzyY3GKQKFZBLuuYfoY2hHPex9ttYAkHAJH
Fk8XLBnT6JFdr9kB5NDiNMl6F1kAgAmPcwkMVE8TwKPwmIMKpYAVALN2I0KKKHmq
pUkfcWC4HtargjckQET1kdNH6/pFDL6gpJ4HFo891ZMd3S4tk1o0WEollyDnuJCg
EvdOPmzkXJV5Ahw5x5R1x8e6euaatU6WbC1xbbbAGb1IY02bxyr8azRGaXem88UM
tIhTE6wPp6FdQ5qSyLWEpE0QZJM57SLgQ9yoMKSfql4ypNPriGNTdDzpetl6qb+R
2vlUh/YC4F76VsvGfli9Mfo0cpH8omp6cH4keraunE1B1yXi+1uY9EiP/yAg8LQV
XgyBdifldh5I5PzpjGYXVUWbDtXyxw7ISt8nFbKcZlurN5nsB8/onJb9Hcc+MKzS
J80Trp7bz6eyoZd4h6WnMf6/2NyTbTocZim2cPHTaFHLvmTCMKl/317fFTth3UKw
COe4PIqOps6d21P+KeZJMKkjtlc8YFFblURmkVpWK+Bwa5in5K1EOl6wCqWU8URg
wIo0qCzqpE7VyYP30YVJpNQpw7vF1dC2AbERj8vb6ITGwvDeLIVnNf6Dd6gdc+yZ
fr4GGQpZog0k7DYer359WDxCM5x7QKQNHkQXNTkOr2QCF5yB3hH99OtiGR6VENi2
IspkPTQkZ/oLYjsL+TAfVcEy4Y9hwasaPbpGDvBjnXr2uKLZHb2/ri7LRiirBPkQ
1sev+/aGccCYZPanAOwJjrg2iw9cLjM9SoYcLeZoQ73TTBFRaIzj1LETGxaxoxfF
5K4OAfh08IX4hxsn3RTIMzYuODRvKjjR/Iija3+rIikHx3PRCGT7TICFkNb6deT6
2dOv5/5e0jrLJiFzvevTg2qhUOqQd73C3jtyC/BSboe+kBfr1G8mo5biPs3NZIM7
IFe2lGVA1qND1NYszsCH90+zPQKouYZoQIGU29STympOEDRz9i+ADWlgx3rux5zG
y4VeO7qdfigRUuoICJztTM+6HWCYg1aDm4oi9s6JOxQJ4XT87Jy/CaEanElbqWsB
x6IU0zabem6cerXDn0q9DmhkIt4fuUKKBg2GpR/STah7pyx4KfefDKywXFFKORxD
4GQE7iBVCjT9Py+LdESNYE5lUkAN5qwm7ui+qxTkECavreI2eHBNpRAM2V6fNMRM
WbKjiDpkSH3p7e5ozlfBZ26+ZrPjWzxO6gXGBfBFkueo3GpBWbkgp2G0rmRSUriB
hwp+p5oR210luc8OoBr+vOZCrid/QuztbybDCIA55Z0qcp8ukE1llNYuy78mbPO4
ToULMtz6/AQC6R53qzTJbdq72lwvGueArp/yNHPRs20sYlQldINKW7STHWWbTYZq
bdAovUOzNh+baiFSp8sJgJAhsGf0jQMW6dzFEux27+W6AZkAt2Yl9WjYsd+MlpZ3
83F73A6i1H5N9arzI5QK5z7CmxZcVuBsWlVTNM39HwoTNyFmSIH+92lVog3634ig
90vvoELH2GTGhR38pPpeFatiq8MDeVn3Xja1w+ZL/uagN5IKOh3vEu02dPTT4nvV
LqiUu5eM6CL800ErY6vVcubcUUQKACakrbfOFZ5GCRjoAsuhemH9YwQoXBkYAfQA
3MgYY6euBwUwXiBrE2YidD1PzDAE4326rAmOcTbOxzgokB5pbM0mi5YdauNuivTL
z7dQm8kBtilgpruaBQ0r1lBsBs0hKKboIVm2ljLBJC+w/BwRVClqdljaHDaWA9pI
/sT8Nx0+Ob9U9jSTIREfGkRJOqIB0TgN7h4LHgSVwnDrMR2SarN4AHIORKYtYabz
ZhS2QoY70K3SiDl0kLCz24qAdomLoK/MRSO7U0/822RUEXgIzHsVxG6AyV4ClYti
08Dq17EgsNI/rmJIYX8EWPlrA4TfJHnjWmlmnS3/uXfz1LH18PMh9PlSbncBKKBK
myjeSHD5Lc67Qot/a0XNGMnhthd1lq7alE98SKUtHKdufbbogmW7Qds4LzsI50Ch
Hp7OtjJM7JyK9J0S4wFYiZGFTKqNnOCLkdV2cecxLJI399hKqL1Fks+63RwMU8Yq
psift74jGRd9y0/zCA94LTdzh4h7nuTOLhV2Ix37FrNLAWI+g3m3ToqnmD3oHbUC
SkmfduxpJYu+YViCoG5w+Z+znQr4ZRujYq93YX4wJBUdhOANeOd3E6MZPcBZ3akY
tlRrAR0hXdTJErFXxy1sJ8T8d4nlTKek1UdvTNgjfMy+rCZ/kAW1faKvFpux1kWC
4zu1ELNEFLc4ZLHU+92ACEUCpfRfnccZpKhHyOjMW7EfErUf13j2vMdQfMRNtKcJ
JVYdzKEeFUtkY5O+Cmqe92TSrNKh3IStEN1h6+dX1CdTHhPGSlqm4pq6EDT77+PE
xXDsEU5mKaFMJ5i8pe6qLNCfFdUmnm2tXb5emADQoxLcpNzxLbqKt+eypasBAuUU
0F3wPg8/ZK0wQ/n8wtapLyRzPlihBV1oWDzCad+Dpk+W8pWdTiFsg+ZIVHD4zGT8
0xt9u+sK7Mj1miZGmBFP5Weepgaa9o++dziiKxBwT3smF8EinLb3NGJPOk3dBhNa
4paKV/nH5UkZcOVVZY5YEizjEDzP9IMeG+fIK3qCcYmES6mAuyDZLEUDStehE+mq
FmgGP+nusm6M2YDcAUDkC1Nvhfj6Rf+VEv2/IWS3MKzFIpMvhhJpPXWZaGQR7Eip
+ZacY05ohmcxUm962CPn4vkKCwVLQZ3JixMRJOwI3lH4oRkG7/9vvZ7WD3y5RfL6
w9jtLPxxVXZyDLBE4xecw1OgQWAw5sCQZyHL1SwRIRmcpr/XqvHY5Z2Q9waobuB9
5A3zlX8BpzPoHTZ5knFXNXZfA4mk0yswCkISDaH07IrzaNZR+MjZQiDkes1Fg2rU
gFDIO4T5sUxLF6GiNYW+kyuiqc6qI4/U1AduxgY3N4YpHvV9K49rYm1Eg6dMp6x2
qfVBd5ak4Jam5XQh8/JsZaCdaueJHJGmj7Qee2e85gRY8udTI+Z/01XUuyAdI83V
ZKZPdfMd+otIsr0gfENpSa5ZlTmq7g7ErTRXmcv2l08=
`pragma protect end_protected
