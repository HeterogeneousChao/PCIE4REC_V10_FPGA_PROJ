// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:15 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lTI6j5sYeVITdLwPVSyQJ8A9ZqMxIQ9d5bqjYdfSgQ8fdoAxJRxWI1cb8Ni4iHlP
6TdtLp3pXjRWSWhVsH9ILLvA4B7gnHrkO+bS8q5yF+J4E4r3Ine9JMQgLw07pa32
BZhmbjEoi+n1JNsPKugjHHQuh848Uyk1k5ldRbbUj1g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19632)
u5hxdkqnmiy8BDoMsFL9iVlZ1uS3vksTfgRNjs0DLFMdwPMQaau1GH1a0tLL+HQ3
5DB1SI1Emd+LC889+LlH/JuTA/STm+i9qGl2cz4L4bBXh2BIe6Lsz9QwKWQmZlm+
kpyYdwdD+Hy6UCrZNwCiTHm9DS6lZ2JAFx5NunUenms46ahSW4ezJgbwzqkt85JI
dKa0QPWshZCZxLMd+ajQ+Oxt1Y5v7wClWaUHsTeN4nk4eXCtZfwRhEAzSUOpUtVB
3F11tI5+TB17Lyj52Jk/9nd7Qy4YCdDnWRJoJMkzDRWxC/yomldALGOiS8GD6cPQ
bQ5KI2p5x3xLmvIyNxOtnpYtcuvenL7u0VQG35O23T+wYoddywPCxsnc0x/T1nDw
ni6w592mNRxUEG430b0XrnthhLQu82nNnzL4Cfb5sVoYeYgWANyMY7/Xiqxpnd8Y
29ZGukXynJwasOrYbpQqqVK/OeOuF+pZHoleMEJz7vUATGRyzi1I/Mnb5UJWuJ5N
rnZfPsbSusdO+A81b4p4La6cnFtcITj67BZ/W3cBe8QOk1FraNnVH96ZGFA5H+CU
ujdjtW/Le4pf4e6yZ+OMLG+aBnfAq3yJWHZWMirojySnmmmkWUYBffmJMmi0Yzhr
KXzLc6TCKe8ZqXmMXzGqk40d1JuryhHwFQup9Y4iD/lXLhgD8xfo6r78JDWP243A
HZIvvue5Jj6ItdXd/fbGAqBdKHwmTOcN76ULmyviIXrusKIQi/ph+jFnXNth4cym
DHff7682MGQAqD3EqPYCLGI/RVdv6fUBNwifeqILmO1BrIXdK8/s9CUaP0MCgNRV
OcmfbrVgbvSPOMwiubzMc2U0BbWVWvBbA1lx5GtDcAK9WWzR4I1AT0inijgZV/4m
s2pvVF+HqszwABSdAY7yz3sO1IMbYy6Zd3CCeljNBZMeyXGAoeOTYAvec3GB1ygP
OdV6pOuesFO7ZvWMj+7Tlx8yOLFI+xYkybWh+A2zFjbRmotKmDb5qrOd7hddlS1Z
+GjlHBFpB77s0srdMywmbJ3lkV73AGUlOifLn7ZEDqS7U7QDh/mvEhLJqD11ssoq
yaEuqyoJUXA6wmgnDjCXugG/6huKi4OddFJajHwdMm5nqG5/JC/4JmdKhu7PP8xH
xphxtCnHV1Lven+veyq8f0H0cY0RYL2MYQvKNl1Fg9s8OpmYC8UO1F34ucinR1C5
DUEhSrRSKkUy9wf8HYGzXmjZKf6smLqmprmAo0M7Sq9WjuceXycqVbQP6a9OpiEQ
2x+fqY96N2let9qkZv7If6IfLjRcmJM4o6M8WaF8O3wc551hmRC66C+xd5sknZtt
CLugjoUM1Eqzj6lX5mZWx1tLIyZnLjXJjS1SZSZavXq0lmqtlQXrIEeO7d7Qgm2o
n2ITuK9yKXBHs4KXUCCdbeaM31v5yovTvLzfgx2qljkklIWrUMBocDC+3iHneB77
66PJXE1UXqEiX+Rb1DrgZ9dPWmkr7pq6QeGII2d7VXdI98mthCjmcQLaHwsOAUoW
zRP0lSNtqcdWCXrvEOVGbUYziHv0jnxFnrKT2t6O2etDNOIP4hICzxJQ0oSGwdtG
v2LbhGa/huMvmw36KFL9A8Ok78J2AsnGCvX3EtAw2b2U8dtbjnzdDBt/rx37UsGF
Rz6Vdoz1jI81hGJNp0YWmYpNeNqWORIvDUakF7IuKL368fKkdeqpd6sQhdrdFXUk
vZyDJZRJ/VvLd5FKOYe/rfHe6O/MuoqLr96FaZ3AIyNS1oL7WLof5BHzyiDighfe
O4Wcs+rbOllydUtq5cqnZIs8JHv8bQRTzOd7tE3gPQyK0Go13sZj/QaJ/cR+8Dnz
pr8I7Ts0tp3210/s8ncbY97XTpJNg9j94dL1I3tmwddEmvWgFVpnkT8kRwdRDv9v
jYtgELcRpj47Dq6580A49UIHescFL0Qyap6BULdHwWNj2IWgT7TLyBUuU4bxZCIx
7HigfP4L2H/7SD81heVirny93fVaGNLOJuHtae5JtzdfRdmlwOYYSmxzsAQNzOY4
pfcwmuJom8BKnUsqSPlBdvP30pYopKKhIKJ5DTo9ewkWhPMDaS5hEBR44PQvUGr7
sK46ztZqxyeR1MxBpt9RA6iFBpYea9+Xk8VqBNncLeGwt2oQxxF7cKMoo4Y98wt0
ozU2qcjcx3BOv7lkZBhVspnmydNwm1TRvNVOMVyXcAWj1EqjwUU7N6W7vnl4ElUr
2RDl75A6fkhypt4Qu0FiyhTrbPqFMyCqu5wQmTXbz7Pk2WBh4Pqrs84RVxnQyYXq
ZnJ8LRu08ssPxsPZk1scdtfFShHWM9bUpCXHkpmfSiR80VDS7fb/6ylYtFbY47WN
tr8sbIpMkrj97YEtftasrCaAqsDg9HO/62beeWGe/4DdWGPk43ifQHB7SExFloN2
8jCoDA3Xr1P2R+Wi0VbTFGkLdXIYeDFSdC+It2TgQ4LvxRD01j3xflagQ9xia7eT
42DzxX3R0ZMltdXqGnlM72jLK2tVpmEl+15Zfoi9rsgGzp6TgxEAS6cRfoucMObb
N17hE4siSN2GpVLID3LNShjpFzME9PDMQXqd8Z5H0KVUcNv1u9LHNqhpko8bYDY6
1jmw1L//RMxKDDfYFywvX7WFaSkjELpDGPnSiVNczwzO2fcXKsMAYD7UWzzDaav5
5v/uM5xnQA/YJoTAfY/5CVCmy+NGW5nbdf+MJpPuDeBnvB8ZoVUccexKTe1f+V0f
E2J/NS7jLd7OJcLHBnE2GtKXXIfmjT/Ay2UT34BKvVvRjy99tLZYhYs45JaOUh8o
zhs8dG0s4eD6RbozDy5hTZIsg8dLJ3XBI1fIazjqsZFjk+UwufTUCcaufHV6NA1X
cVd8s2Gjs2g6KKm6mPdvDTS8Q57L6UabJ99WiXanmalHQcTvPlnf/q6j/M4GUlff
YSsRcQijGaXetLSo76U6E3z+8EB9/LV4l4Q3erNepUE6yXKeKeK9Orwk0meGO4G4
ily168xu+yLUl4dX6HO5qWRSp0cZslBpoDxkznNw3W7mzlwXQsXGMc6qCSRFhrMl
6SBpbOjFpKW5epTkB0YFbWjxF9SQGvw1Edz53fA6QrD4+cFRPz/gwSPZWxkKmLTC
qKPrZmMlsnvixET45/r7RKVtPLBbj7b2CP2Hevd/UEYQT9/3GW5OnkpDL1LMJYij
Fry6MxieGXr4TX4GYGIAaHjx8fr9f1vniDsfylS1BoDLVh2zsABGWadunrEpAEcU
d1FktgxGaZp1ILCQD6T8D0R+FVoPO9ZselqYLnpMRYxs84CsTQocggKMW478/WCh
p8SHgK90nw0u8c0L2pC6m8Mbe/wpvNCIJzW8feERUPOQ6g0QL/+HarRPD+W3toTy
GfOrGnDmP4Cu+vuqjIn/DI4635hxGTiWp2/iaKrH2hEKjX5t1xIERJc1ozuk+ZC3
QkE/kBBltomk1XUmoVifFVr/OIP8uhcqoskbNhgJw4lhdORZ6acObvB0NuYazopd
96hCjC+dl9/uAU7twy4Gb0w9aPxW8XjdddEM+v/eXfUv6IRqK92u4u3Hdm6mTUq2
xa6naCWYpfTgy2ldmCHJNuxWLXJgvi4hvmLC1Fk//cszVe//a8h1xCk3Q40Bwhhj
Cj/2AZQ+Dfl+ciOR/dUiApOSBwu8xFnC15qF420A8ho9+zNhwfdi+DRkBU+eE6l/
qyTslqM33w5VKDVc99wACQDowO8Ni+MKkxPsw0D2av1wpEHJehMpT0XKqDiODBhb
hwDDtmLdEJu+Tase3EqwIIKdYt8t2uIpYKpXAq2Or7xYLOb4zfJqfgTDrQv9oc0J
PdvsrZWGrm/qy272mtlUnH0SDKpBPvpLklz8Zp2O5+u576ODHW1+h/gUfP0/w9Su
s/1ZFR5jDy9nd7LNNmfqHXobd1bawW/Dx0jokTWEiKP0OYSCUoT3U56Pe+i2YAK3
DkPsyp+FOKniyj2wiePm8STr2mLKYfQDwG1UK9uVTHU6fa3xVaRi4HSR1EwJ2a+P
bruueIfLirFLJDgsjspEvLawNBb2Bpll5vktr7DmBPSAFmiCPWLMdvkFoOaRP8BC
UGDKAuMXMNchF38AmYnjEqUbD7046tPbO+AuPz8GC+2bCX4Yez1/zuT0MKM6I5BP
IlD0GBpXnvQQW0z1knPVoPNkuCURJxVWfb6RFsP6YsVm5M1glOWLAcrRY+e6HCCL
4u2DkS/5/Rdr8RX5tRW6pL3ByxOI96kdSaJ9ttT6W1HEsNEwPJvyfEgnTlmdS7lQ
EMkTOQXrPsEJUc6qQmzEtt9LCtVKPjWm/k1bu6rOrDraTwxFtfE4x4vggpjp/9M6
Itrm9ASbJjHHfWsQ/H8bdQ6pfgXlnahDIpoSc5Ak6NLZhYlH1YpyGGIFi0fhymT4
iptzCIXlhM6Q3sIpyBqTvU/dMDFPK/jPwLnWoFumYizd7Rq/jIscZBpMvjYI8fkP
USkwW2sq3BONhyGyvvCo1Cl4eEMB5PYJqxy/TZuRjoizxxJgnI5CbJoM5vijk2Gd
cPjLx6Voye8y3OzOiV9Pay5rZuR5UBYaSUWz+0DHJB1pGOokMhU7cYefG414u/F9
3MyNOmTD2pyMfXF9//vyudLLSjCV0ynzXfsP4ZI3QNSrY1ZAkzyQYQSR21NYctpR
0cEZFNkapB4Iuz0p7Ia+G/bPPbJ437X2oh8OlnQnfcRO8j15v7BfLLjh+Ev6mviD
ORt5d54f38I9N1KQ/ngc/f+K0U/zPcFbq+u5guBHWC5QYta/yZponQw2pV95EGD/
KvdKnzisPAdsh0gK90rptCDfJc0y0SxkdA8ha5dlPtGAkL/g0NMJ/A1SOMoHMHr5
rt8ANQdDj0MWXrj21RMx60DnodaT7CXZdz26lBY/qODrsE/hYTgWDWvORNjmeA+b
Hx+unazqrXqdK70Vu0RpZuuzyGq+nFkJ5Ki1U1LgUVr+MJloDQ5OHTSJ/Ym/Ln1N
D8COf/yfTjXd/L8G7qSig8fB/tb9TY5snuB0lX3B1PVvW71hNW5KDRuBaX8n/HEA
gYX4zIbKKG+eVPsgmWme3kog8mLBLfefpL3c2gPTPy5e7Omc8Lq5HrBbUiWHg/VT
Tr+uR1FOcex2LeJUEhtSkaQIG9BYF2ZvPmwni9y8kKvxxKFssqQY4aoNDXMWdRNT
KKq0JCMRfAI8WEBXM7ThDspNMU14dtIBJ74nnfHmWEitoYCDrcUjXa7IoSeFZ1nn
XwQxWIi1qe476Jr3aCO6TNjfQYh5EBM9M66ASaFH+9ZiTq1vW3OacHzaKDlkhlSe
+cSuTL3KAexpf2dQXpkXSh0tCleP7G/HuVYnrt7lOBeETnV0vJwn1NGjDG//lFbh
+AZ5qP0pE3kxb6BQuIomS/ziPjLCCOk83RmcttpNvgAi2TCrItWvSsU6P3em+d8i
Hmmq/ZFZNffpvqg3RBi/Oy4Axtin1MugGJjxuRsvxKehtGWh6JvnV+WQCHpmHBcf
SuMJBRXR2xh855Iz6ZWd4eqKPqvj/riBc2GpnzB0onzHULqgCE54ubW3Ax7Ji2LZ
0ZqBW3yKFKWXzH++KmL/wIxbHg+6zsD0l9TvnmMo1fnVh6MlQn0v3BJtTIL1TROE
lVcwTdZyp9OmVjzjNqpP3d4eF6t7XajCbpJVbm6F2ky0Rse4DSQtf4NCYofBOoBb
tyzbuyqdGpaXHTlSg8twp6UZLhvBl1rPKPPm7LqKzEV3Y/6MxmxF0WCHfGPNeFm3
SOhB1qO4+sQ3EZXTo74RMhDD0cDdRj4c14+YKcYH65QZJ6HeNkXMDxXW67YagJ5O
mL0c8F+4p144Mbc+wzkXWXUOebb1s1Lb1G0Jy8EYcFlP/twGsktg9bwag3iB9tmX
DWUAnz/10lT1saxVDIeaLV5k967biICSc3D2vrB3sqGjDsICyU1A6gc7u98VT+a3
JbP9p8dv8pNEaRLLzFddnCEv0a7UT2w4bI5JhXM7jyxpyg5OR9MTGd/8o/0naxHc
PsfTJeIuShyX1I1hgLAS005c5Del/jUUnVhvYOGnJcGOto8bs1zNBOhRn+DrYVHF
vFeDxeKMwuBbGFmj9ZqLj8SqIXFWPygAtQ7kjzmvGHx7SMieCLGwORfR9Dr8ignr
ai8XBzv/nrd9CMVAjCglFlyAi7x6fZhx1kvYjUwfO/qwF1kVCpZnVNrP/XHxEE9t
hNnKmI9cZHg3sGNEzp3Gq3sqq+YjVIH94kRCtPU3grYUlEl1oIIoHVBRFFkV1GxS
ZIGR4MsckEtUcaT0gGNZa/oKlO7YKq/PFQpPU37u+1BNrJ8WZE20S1Px4CCtJz5m
gRFhZolb2VXZAXB4YN2jhHvQFd+J6vKuRxU4ADCWg9PqKFTeirIC2B5z1mMzaMcG
nxDCItlbnVXcd7snNGFG8kqiztS8uHzOgXLRsHk7TQ6T4A3DicIns+LuZlRwJFtZ
xneYBykqkI87LQtWqOi+Bw96cdS+bNv1w7TruiHjHL40b1wJ7gIOZKnpsOX4hZ2q
Mg5sAxq90mLINSAuv/CkdotjmjDYFUyeNAp1l2ilbe88dM6xCakc6y/YDn13P1t5
N6PNSQuKTV/lA1Uuc9z6EmVeZ2Q3xOZ6rQ99nWcDxJ2pKPWlX7GBTzZ1m1KjbL5Y
vY1jNqazUDoQX4iQrjp77ANXQDstGJCRh/hPCk4TFZ3bgd5eWP0KsQULVWDEp47W
/BMfrtQ/6+z3dXqqV91VI+kM/pErdrpIDcofX8jwE4l85w55eyxojNnAajSd2cZe
6SD4uNgVfvGlcQFPWU2DxY+ADmYHTcWkfI6hEWhfI21FAE+UzrlpKgf8A8J6t/rr
gppRyD3BDN7DwWQcejWRW3V9tIlXrjijyJzktSYVaeq0XVqs3zfUocSs9+b4CZBj
7xxHvwCRRYzSmJg+maAVGBmodBnlb+gTi3x5zqxGAPb3jETcuElqa8J9/YaB2r8S
ZE2sH+wnwCyyAUxkWrZN96bPILCC2gpm7BV1Y05SsP+BYkdwhrzNXPk2LTfiyz37
WLKgyH9P2py+dv6Q9TKcJ+VmRNXX7ssc26tp1cbUzjgsSAYVJb+iHLGxQ+PdAvSA
DaDF8BWoOaJZ98GVH9x/iVV002/qkh8OX75ums5hsGGakewEgk5pW/CeFIcBQYq7
IAxTLeyprDFoYq6d4tsAAzTMxvlGoSqxGoviVHeDybAGnJpVJwumkMlbIgOXbKeJ
13+/1gY442n3n6D29q0F2MsfwxhcKbfl1ReWJGymN2c+ErxMTM0jxWfbshX3jgpg
UsoQStxnFcYKSXS3vL6cf+ugeMbw71n+r1++R1MRKXsM8kjNee/6Z0EkYrQGb/BW
ZKP4jO3JeTkkZ10nhB/F7hNoS0M/yNJTj3hmhw9c13qZ4m8XSp4iJ4mVAGvtylEU
FyA176YKD0mAx8KzjFyoPyfUelsGSOlG2FlsXXGy+wO8ML6suY6CTvDHBNAiy8NE
4HOsErKUUlpCW4x3Ot1xbS8LIvpfvUGajKkYpb2jvtRdMpCtvW+fzPOTj8Xr4Qz/
tFiXAw1jJGejZHx5Mi4Iq97IpwRNH53hlHYyUQVx+8Kz2oHc56tp/DyfsZ35c41m
p3xgKh6xF0ImX6ORbgFNrH5uUlcuVLf64BNvwXjcmbzFw4owfHB58Q+1t1evu7Zr
IlZWZ+vURg7d1F3uKhd4ibrl21Tk6DyIfZXe2mC7yxzUwJCkuuA6XwMpyD88HbQD
kToiuB6uWtWvsRK0wNzrCXbc2Ra8mUp2BbcTMm2mrJGKaPRpEDHAPoH8waLnubX0
A+gT1ZwgmajqbtGx2Ar/cdHrgI7cmkEQUj3IqwtYPezW1xgQFyEBAhFn6trPIqHA
NYI9yHRhyETPgOCXUI5vWbT59pm3awi+vsYDQkiedbL8t8JUhmnrq5yzscub87LH
O771ND16eC0wbcJ4D9ku8WX+RuJj1S+mNI6vmtLqtKPw4tb/HHSMYQiOPDuhF510
07yY9S81v7tGjdvw9sJGNR9ZPh9OxtwuS5bGirUV84mT71QU5tJzywAx3kLIzd7N
mQNmjf0kXLWFiADfn5DnlJEB/vnCXc/y+C8qSsTeQgAO1hS2EG0WXGibmVBHaDBi
Ruxnh2ibJBbUsNeLLRftKb5Gapg0l73zsKsbigYjI8nUTT2M5loFSAx9s7dZaX5k
WYPDFuU5/JRW6vqpRkYqzEN4lCl+Ew60Tull2JHEJjATdYtA6nLlW3NytoNKksH4
+HLMMnOZ8skj423WQeFMYGNfBAZteprenbUe7asUrSfAcAK5mOpS0c16Q/7bmDB1
f0sFFdf+xaNo9EnfIKoBCpiRwdeWttIrivb556tbiei1dCOUX+sHnv2RGprGwrmJ
4CZhSkkCow3oz101B1BCccGjrbZdzx4vsj3kozo2WUn2X8yGZd7E7FEF7GL09aTa
jAA0WhlOk42JTo+8MXdT87KZty0Inrl8Ft8KqMa64Rwr0kG6Y6s79C99rV15f29x
rO4LO8Zta2n+goe5Ul2Dncb3kW9bV6+5hcJHFLlwesbHEcrb6HPet6Y17UBRFouA
my7dk1Dvrnnbl5OVRc+c8aX8yywGcVrih4XQLDtT7WRr1yb9yvU2pSNpFw3hA4PT
9oNphyjfpGwDuFLeuPh+lVXFXfchGi5ZGhxzXFZh2Rf9sKdIoBaFtjuHLsqG1Ou8
p+jcYrNADRs5e29568t8TfQCNclVqMXvrbAdUmkLix+5GsQoJ3n094Wp1sSax64p
bkyh3Blkmh+9sNVrWuYEed1uH2zPl8aviwX7UlZvtYV6r/Dic8rOtjQo3gW8iPlf
ak4IwUy9IBkN1O+41ns+5Ts+XJ9CVdTd1Vn9zDJefTM37zu8y5BbiidFNExZZXAJ
n2CRpCLlDw+rOlIZ2ry3gvtaW9oTQCdNq4nH9qQEqwegYjF/XSkPycXXoEZfJNne
3RpGIrutKXkTT+1v/h4bujAYb2cy8e4O9NejzDxyNfsQimwx/JBhFOfWzLLOOnPz
6jPRfvx0ajK39pzXdED2vV9VpGe54YRfP8sZjC8y3MvgTTiBU/hPtMEvadp/V9P8
GBEyDwbGjoJeWBY12YUKyIWV5W+sIrZDQM3sH6qTJTPBBxAnrTGKmXJrzVys3IGx
r9aYH/qi8pcxe87mO6re70qthqs6b9CaTD911anDpKX5jwvIuGfny7T7XVV+wDCz
aBctdrYD0mGCCxzNOWfN0uXEkY3+UUuiI+/PQJPHWNxicAALKFLDRm0SXOO9oPe9
kYe21nLfPuNC67OVr8MWJbWRs5eWMYthAhAL6dWmYF8wHrpLku9RhvAKc6Uwz4iv
LcoGNXMt2FPiYo1Y1CYgXdnB+5avVsHxUCjK+6gYb9w7QAPLeK9I5OVA4o8SfIHa
LeXyM8+zuCSByy4jImiNxrXmUwsAC0l6MWIJpLMjUHS8dzUa0NxCuPKsjsOd4ksI
fDlPJ0m6uuvkkGPADW1V3k5151thswAFOepj3refLZW5Hkg4OEieVsagZQEXfO8z
xSHqgPXmXUgDnbJMOXwj3qFTJzeWyehot8+5i73LcQnYH6fPQpaea2ojzKYxIBSl
CMLY0WXN9/9v7Y1+fWh1jP3e3WRHeOfZ8EaxrDMFIEPIZl0Uz9U+9q8Ev8805yI1
j7abJDgyhW4udzdhD1TTybTFh05XFQxdJRDg+hZpBtPlCC8AT1xKioL5qogoyzlC
oxIZ8spK6NbfJO9AfSSSqexQC9WNt7vZlKr8AJg2ThJ7GzUB7NcbErVh8IJvYqCm
hm5cfmqDxoIsHEVwvnDluoIiqZaVy/wFSvNpqCpz4v6XS14sbhSrHfIsyiLaZV8D
gJ7sjL8ZRM/BbsDkCRYRv86bRF7qv6UYN1uGqAIHb2kw4kuDsnrS3PieMwi/LYsL
HWqLNLbzlFGce5EmzXTQr7fhMx0FrrAskdrAc7oYMqIoJRnyZkafvDz3haD5QiJg
Cp9fujton0Ku8cNXHK0tWSVa7XgrNdyxz3DmCheB9O2K/JJ3Z5bZil43qL/Cr5dV
XfHv+YRGyNqBV20UkJwi1f2UyJOKsYb4CcoazsyjoABOxMI4jnZcdff8f9k19kCk
7feKy5OKuux7foDpv/YZbfMJxDS2cWZetZdKqu+l8YV6Rqytj6oKU6Ak7aOotSIM
/eUxvLV+JSDU1gzeIdjyVKnnoWtk2kZTJavs5WHqt2tRCM4ZwO5K3p1g3k5sUbQJ
W34Ye/3CSHM5plzTIBbnbjioRRmLRV28Z5DO/MUIlFdmSYwyJLgv8fMIJC98godj
PS5h4H3RlYjS18HTJt09vCVG+sKrg1eoglwdVAv48n/dWl3uxfc+CaKaagrjweyv
ZwB/6GHJXxSxZ/Y8xyO2uEe2Ado0Ji95Pvn+F9fRxtwD7JCPkVwqze5waH9PksOb
O4l9KOV+Eylyp4XyPU1nUm2IFUYF7Mrntsx7431WnvOXbg3XQr1w2tjJY6LQ++qz
df9L1xqDM7WALQ71KJJ4veMHl+DOmgd3fxgBWye7yqwl8u7cqfZJojmFAuvhinlU
1inN2arM8degthW3AjtMgJMy+O8qAdcMQOy3XvXo+nMx5yyi7SEZs23fO8um2o3l
Ah8HGCf3zZP24iwzvCluQ74lczgkHEw3vhi2ImCpCOXi94E4RHBpdOsgs+g8Qb/f
G/Dy+0TM/yGmDSIC4o8gWd4uaoBbMlj08WCqNYD3CHO0EE1hjzObicv/lj92yjOK
x2w01ehwpBKSPNjcB1ZmfEg8le9RDM1bY89w1S7eYcYe2i9WeyGRj5k5JOOtolyN
PecRvq/R3PCZ9ZVyafNaoqQyYbnd/xCxQwVeFvanKbxY4uSNKT2kX5KPxb8ZoWEN
nzqxuthnkAJX1fG1KooEmWgB9rT4gdaidRlNT2B1rbcykmp0lPt7U73tSPEJ4oHW
XazJRKIJyQRUtDmouyo8cdVPrwMxzekL5bW8OKDLuzLUiECPn4qBZq0G0zAa4s31
A4QB2Y+G7guYZ0AH8adYgu8iphPwGPoczvYlExXjgErqQTRu252bs6FBvRPGlqgV
Hu/J3lJ4CGThLiNzWkgthRtYPeG5KiSOdSRntgUXxYJdqo0hstqusb7e/7whHPt4
RWwPedFyuXU60/WJcoV9Up8sAOBu64IJQHVGYXQuOoL2Liw/UfxN8nBNZfLZygLv
EcgxJ+MPrhHvUBXoSqSVO5u2YtTWFBkURhjzj5KvKLFkhH8g0/NeuRyj0H8jdLdb
p/9kTG1ESWkrFApiQGESQr3xwS2ro8plt5XWxdkiLvYos4b0Y6Rh6qmwXjPsXD8H
+a/p4/IpL4m+4ytR/AXgnIkqvx2aqi12EOyn4O7AbPni4Q772M2mRkCCCYCT1uLS
1B9mQmWtgXMJBsEAWltC0PYqkW5BnA+5NojtCYPPXgr8GI4zuzedwuZkHbbRMKbF
U9WAaOs+n0av8nVbD6L0CepUmenM49eeoOlae2ojIieddXl2THeLOwVIw+8yeC0f
HH+O7w0ZZBAgWyfP3apSoc/KOUczGJ21jEnUBeP7yWuA28eAmq/12wBvy6cbGLGv
9sJR+LWaCsVXZiFBxmMGfJwJawU2FFCe7lLHZMLNHKePIiqVyUkYOPCxhAZR4rDt
9CWlNpKdwlwLd3Q+nWEwqpLg52Vk+a3p2UjYJuz0Roi1Q2E5eJQmVWea9BFkANTe
j9YIyi8Y2xDQtMpiwya0L2Vlx+BpgvFFQP0GmKXzHs4sIbGTm2pO2EdAlWbC0ojE
jkyf4k2YJrTrYK1oTVvqEBoVHK1M77MfA+op/hMMuX/K1A77KugwpW3wrjasJX6p
uRsV4suVOWBdxBojNu+xPbdbsrhGptMHD9bg0RiPAE/W2hG7fg4GJAJLIrGYKCfq
qCiy7nrjVKYKAE9VMpuS1Qy9LkmlW3F0gGaJYLwJpy83FIBj5ZZEpbokzvK7d9pv
+ophhivfMV1pDv3VTr0t0f7z6PTDaYqV8oAqsK9I2HTgdpebGMs2LIA/R2mPh75U
l8vNxd0DEsj2C6E1WpI0xMHVi5pQ8iwgPHgkrYeaIqsJCsvNA/sHBv8NvW3sVRou
T4HoMwwBqv8QTBCTf8YAYDhZBw3lfUJzdrM4y25VBrhkevzkaTuRUPQFkNrlbL0h
Kx6ZyyYMvBgvCaSKnltjklTNOdA0ahRbjdRJ1HHpdvPwFNqDIsv0ZcABPUCWkBHg
0FzYyW921KSdMvozBksz9Y1hN4vAeS7e/Kj6tMA7Yq3YsoxyWeyom1xUycozR7Pm
4a05+rCYEUhuKt1Lr0OY5QIpYjhvt+Bk9Inw1TYKkuHXxv6ZYubtJ8sdwcW5jtud
rpA5SLsXKv3MhZrqE2fFx0HrKS3zTzxNsrLk9VRneLbEjct+c2KS5fwEe1g1aArK
H3CfxA/EZOMaIhuWaScgBG/gCw4vP7Sp29av2szuhB03xFKWq3ImPxbNI+O7i1Ti
6z3Ugj/jUTwLBhkA+GMgazPBggDX/KKhzf5B9Sq3SEm2a8/IPzmIXv4vG907c/PE
/J2WqYoEO1YkHjkpWldrAUNbe4iVXyvJRmuQRcP1laXnI8d5LW5cb96RbeUrvBsN
kwcT/lgFAO7eDkg3LL38jAywbVRNdzh4NJuswTt7fMcCxqc6miRsSSnpBP44vL4V
RsnWOjzIJ9ZI03d5XHo9M1bKOcDaGTw3mu6TwRN/n8VG/O8P/Q+uTnEwv+tlJ4Zm
v3Y8VTx4jQ528MxfYFzwuTMlZhiuRhmMloVC54ZOB4GMc2upzU1b7ZkTGXt+tFu8
rO8YZSY7hL1E1u8tcwNBpfZ7Sf4ys32ELQbdLcndm2aRIm1O3RsyidRGUEe7Hs8d
typ8Xh2xjZuAcXUQt0apes+g3yrGsH66XuIVmQUJH4MUzuHDQ9ZBqiRqZBOcpcfE
i1VaAbCh31HxHAPJKX8zmhFqC521H03NvOTXExM/ChDrtamkHlk+4y0ynGI4Cglj
IR0o3rLFq3m9qG1L+eREVvm5nLywXcoSDRaFKWFu2dWVu2U5ZMHMEp7MPA8fOCzO
HL+KmTbAzOiwfQ2guP6DW2OImPKOYFVscTwKJifGFTf+x4LzgbzD2HB9wrkenRLj
W/bsL4JH1q6ZEHoEXfO4KKa47fetHOWAI+xD5upFtSow7PdZFuHv350exXhMKv8j
YiLXYsuGqj3zxYrdpdYcrppJQzSVKhJ+yyF0jy/qPy0r1cdTxFga8F0aZ45WQYbS
IdNfwfRFrLvTicJ1+dV9J065cvTF6skX/PiCGH7ZE6boEc0GD6iykRIoc9WKavHJ
yeRTDROpO6sQI+fI/Mq4cFr6Pg9QnzXjToKZaXOZ3vLMP7+aXTRCGnsKj6vAKwv6
hE+If/l6wT7yw6sJ71DAbbzhN7dvuSG00ebloTS1Qy+upwkind+kafmo/+CvKrTq
yBLl7zh1Iq2EMKY7nNGyJDuFt7aBA9Dup13wwvT0yTVFaI394NTdgNDxnClDwfW3
jBGimHWIpy4ZSHkuBKiDWu9phUeVSMvrpQPUp3FahCcHxDuR1YyTQlLq1lqorrM7
7Dgk3tDsMt+B8Ig7TCNH2OZ52nARKnTt6FuWZhTot/bzOPH+rUoHNb4mqEeF9P2W
/d+S6+tmgM8EcMrnH8nQ3r+El5aDn3K396b5DN7aP23n/TqZDMfZMSUkQM52UutL
NvFFXlNvmnsdMd/CMMnad5NIGKypLt109Feo9AgrS6QSurFs39njINuTZvC6xWVc
gUEzjihN4BEAgVqCda0Vt1xpLQ2cci91bIyza4cdMEnXLDgNOMDYVSct/Gf20D7D
rBGDmjWiFCHXZZVjIXvLHzL8OozWm9GtaGGxymgMWv7txeh/b3/OpwqDI29Jvb2e
4CKWcS1ezezRQN/apSg9CH3jCbjd7v25JHrCuQShv1GaKtvlW4QVXdGDeYdYAeSG
Icrx1s+CYGKnDPrDCsdD6ENiJR/Bj6XtdIjzLre+U7KLDsPB9RWoLBtrqsc2WAYW
EY7Ex7hhAZJpz073W3vNYRZE4zqJn/bw8wLo+FtCislE8F3mhcGZ5yqxoeoNHd8B
EbW0f7qFNUvytDEn026uQdHJ9IJWZ6jZe2ysZsg9BRlgp5M1jTrmIZLzFUaIggUY
fxW485yge+GmaiPseE2To9AwWCb2j1V1X+qUPCdAfC4R5fhRhKifI8oTYGZ2nFsq
04kVoQpnRBLsYGIDDQgNHJWYLyZHfZBekbBvFVfQACiiJFJ4bm1UUxhMoyl8gpxJ
J+abvwkAETFhqrTYuRVisogR2RCA+CGpQWyRFRlvR7xkvPddEIWmUKggvb5y4FPg
PCmxQIj3woV+1zDv9YOQ0Y/IXQbZui2I1o4PCCbUksJsNdzyxcyIGL8be2iA3Rj1
Fu1mziaOX/SQHwy0nTajpwrZP01a8P7nmc+CoiW03PhK45kr02zTMaMP0D5ZO3j7
kfJkz7ALir6CW9Z/delpz/4Y6GVeRkeh9cvWzB+FW3Iv5h7UO+N7E5XGTbTWb9D/
ewsGT211Yao/TcUXoGTmwe1e2HTpB8mQxI1ML1cKcDZyQaDm0Jo8v8sUam0fjXxi
HCejJZDdu+9N1u9VFly2OygiVv7iPUAcimo8EO3u0FWc2uofJgLz1JdYffbfqUDA
WrNzw293C6P3UtxeDi0k9/VrLSWiDGFgbuqaLYbmHKE21bFQMzd4/n1bQ+OvzEIl
3puOdvM7PMqCnMCayFrRcmCiSo4b+Y2BFeqPNPvbdWe0z0lCcoBbSKUDDJf0vUVO
Ck5SGlgduJ62poxnoO9zkm2pJH5F6RhWQcz+u6qs0dSpcdze+ViyXW7ie6AewjNp
2MC3OA0O1x9O45rFkqepjAHbxhEv+pf0i7AYRWCMVMug/TNyOk7IBeRoZGT0j9sK
FulfEBSRNoSl2Jutboa5MOF2vZGNb6LAR+RuZGWoBNuSfqOrXKj7GrP0sQtfmKIA
uCkDqVbCTtgrhpf151Lb52HfmrfAK6tFhp5efZfTlOD9PVyQ4fRzznGYP91Y6NeY
pmvn7rnA46rQ+0XIsvd+j1tpvTAHRehBeKU7w9iAw/bnY2s/f15IN1s+nkTDeiLh
nxVC5ZS7x+32fGV/HK5BtaCX5sSp30HQlcImJDqR/e7GxnTsJDthm0cc2KETGbD1
OP5/8JC3BUhVlGCSR47erGAj51cxDRgT7HH8eJrPeair7wUF0W35CHuMah7ZFlfp
f3X8l/jQ/RoXToitRgQ4QeIIPxjxvH0IiaAAbNyihtou4D98T2K6PuC89noFAqZN
Z5S7kgKXQXxw+enfGrYQ0MDXUr38k1MIJGT6nxrh3+vTNvJbb6P1Ry3qvZsoEY8F
ph7RxvtwagQsbscTjozT2bytWP0L8a3+bfHpCzGHC7yhogGu4vIhpw7ZrpuW1o41
UzCIlO6SQGJkqDAFE42I45fyruDX7FhGqHX4+HIPVCsa08ew750Ex911GY6XNmi+
iiQMF8ZtJub/LzaeyKoHTui3uIIoHxGJHK90Qb7FJg/MCXLZHR4Djqmi6s8QBanf
aXHwLyL38AZsGFZtaf5ywJIOgubENUSWMu20UTMaJSOdFt9SU3E3EZH6tYN4zKre
h57QkjBPqPesHy/odou+ppgWPehDdoT62Espn+da8ZmyKw6dtC5z6rpi2xt6nhdq
yhgMNjnuLNNO7t0A6W+7Ur/5HyU1D8lsbVWVxB8F18t9PYVnPis9AnrHWjnwBIz0
jDJhnW0gn8eGqC1CwihRWmoqABfwcdYfZ51scjrMg/KhZTvLbLUP8BaPDgP5IQ6h
0AwZgOasoty0FMI9r14c5jAbU/NITBs0M7fzGss4QgtRudrLRZHNXZKV7XYoI6+L
ZaXLkmNP2UkVMoIwL/L2X3NsI0efJZGPdPPKYsrwTDUQBHtNCXf5VGF562q83fa7
SVXClH8c+WEwf6Ek3viKkiUAZfIDdwvz3h5VU7oXoyflod+BiLbAsN97QlVaRFjv
ILNKdkWebRTH02qG5zbcHaasgfr5tSNKsErZXhuq37NGFr3r0/+pc5zgMLSpg+Jz
ohCXPu38ivTyvV+bCRt7E2CSOiA/BO1QiXyXvV+SrHfpGLQjEJZGMFgwOpZhVGyZ
gjqTwtaBXPG6MmWQHJB9klDjqPxB/YgDrb+2JZGQSB/0pkNQmCdPW2BdTbmZTfnv
GmuaDORDD7OCpzjzhVEtQuTn6ctLdHPFRNtFlQsZokGpnvoje6kFjlKKQ3WTemgC
2CsAaeK7d5Om7vtJ2hyS3bFOEPuTzGR8VuHqlhpDQLbIkKvLvQe8yfIpOJNUfGxE
nnAKBpvCKRvyu5GXKggM1GvARAYK59pLjJxaCb0t5GSeZMCm0KdGZaOhzfXVwnQZ
3Dx2oRh7KOzeFPTs/Cykphm/Aevj9UL8PcSHtJl623GX4dvVRrLV8mAdXICaAHmz
f8pcyeL50MTMPoQKKDzeV3AajBgc8IRI09H61Kzwd0If//++3jprK+1Ln+C3lgiS
i4GffUn1jP200sFrezMRSheLgwoq9Dzu/exwj6cmURw7NKiOgQiZx37LtBktO8dH
wtw/IGAbFAy+LITWObYaX29NLsTnbclgxHLrwNRK4ktU+BJk5MlJXG7uV1jZwdOf
tuazIkPxb1Wyl6yyaCiEDWUYVIb8heeep3GsjFbnmmwgKFs3UXeqDUKydG61nNZC
sL1Z2IlhB8Fc0/rejbTYQRDjQfxEt7txymqvQRfJTRLLtiSzY4OfoiHyESAbs3u3
PFvunnF/aZrRynlB9nGQ08n7SPjpOjp8OJSQFge1129w2zo+XpDm1lQLgW9EQerN
dpL/+RkupbbiJHO2a8zj1yicVz0MPetfUyN78XR1R6OY1ODNM7KCIdEtqkZsmxUQ
4iF5w/nu8R3ce6LbAYFjIjUNkjQEFRi7Zlkoo5bnREoBP1a5xMqxJJdbAT9BD1R6
CGymNUeAG2lF1auVW1vdC5jDreVUdc5rPq3YOo7cVOlgtsk/g48l88jhX24wlg3m
AnafuCvof3i5eIJQa2otIvemxBzjfC0kPpHPGrDs7suiER81ibPInK1TeDMPp2Bh
H2xVdpurD1Ky7Tdyxwyvlpd7Pe4i5yYatnVDOA+8AnsaFhHjvBQy3dWImom+54dg
C1uU5FVKyg979eNwDwwMTnXOfCtFfM7LWij2PVgJa7QvmtraLkHKj+ygePIrnG2+
6SsUpnRQ05ullyl38op8+YLm72mHNnmdChDDDpqmhM1V9h/BGpByahjeSiLfF8Ec
lM8kgBWwn6gFIlRGo1c4BVHjwr5adrzKqNrKxcRuHF5SObA4ToXErYwCTzdmdz/z
41Jxror+rlRvYG2WTOWoCLMNTMI3rDfEMJfxcDDHB4f5tz6sz3lHP1/vLAJH52CW
lfWu38EWGv0VHuFcObH9Ahy8YSt/o7QSJatvCNL8icQ/ocXHH/24PDNEhoUn14tq
YXIHhzVqmjq+WY6GWI9BsoqBP5yI9X/75ueaQS2LrSLyKsutX5qlfgVTFALIr/0h
Rh5f+bwFZjYpvARqlMmoio/bcs3i5TxV6dnl952u9AGhaPzl1HK7k30wg3NOR3Co
ugXBsE0U9AOoUmXi/ulfSSsd3gTDNvTfTn6/KPk6W92hxMpaioGfO7KxvCrOBD8S
SABlU7tw3tVCaL7PtnWTxlKQ3PGy6fO5M/Bi6b7ac6bzzz7v7/l9AXEPbvvKYVji
jjta/yQ1jQCZPXaLM4g9yXLy1ee6OZO5DBbvbY3Nc3anqCWEirwmEoWbQtIyjwNx
u5g2pjfiubhnpjnaysp8QWS0IhW02Wdl4Tb9o0/nRS14YGXTjzFGcKZ8tSdlCSmy
RxjLQwUh/kJKNHCFzGwTrGtaj2N+7D1WIWwJBr/PgkeSsi7vmYHzEAvWPcV4ItUj
z5eoAv5MM5QFYkJ4n3zAU3cNV8KIUqrZW7+kKC77MKofnXlCKwyBWhODAkea31mA
evtFOI7Bgc308oRIYoRC3gYVpOJhGrNFKLCJJ0RmV/EOzR2+vy8RZ1PQhVMYC/+9
Q5Kjn+hB528GzW4vPE7RSVQ+3w+8WvORfNQUkSmxivTEmvK0wxS3BiXMnNA2iqcx
LFpoxMfy5MtRYdRmnNScTEzSZtHiiry8z0pAPGythbC8HCt/P+95w+hQG79UdJRJ
5whXB51nUQuD6dv5rysirN91aQHc6miQSvBxVlZGi+Xr8BZAcW4C34QFFZYkrSqJ
i/iyyWp+hCv6iQS5B/RNKq8H6p4NDmJAuMXa+X6EgeDF2dGQ2XFAZTt+k++LdLkO
R3F8dp6YAzlgvt+4KE+o/WvJvt34oNi0G5H32l3jJB/X+8EV2WLR+KdH/eUxP1XL
RYUBeR1N/rSekgn+GCyo6exoIZdVZ+ptwnf6gRKFlP0LnzNCvUkuiQGh9oZnhcwY
mcdeeiHMlpkNLOG2Q7DyKWBWRYalEebJGjPZoAhPxXAV4pKHpmOjPopVpzkQyujl
1mGjTcqpRThahBZrOZJf3QCcUV/BWO55mld5Xe3u/tD4Q4Eoj5mg6ggydF+9JQfO
IUpHJOy/KeLzPMax3S6K/rzcLHmNZcw7C77s1qCrN9T9wjhNlL/tsakTW8T3+dJc
ugQc1RFk3blF8VPBaSe+bMoZ0xqvPTN7H8/ePUfhnrq2IoU+EP0Wgj46IU1APTSm
ghZy2fhXP9XxwiB1fI9S0969bDW0tYXSZtaFM7T7xgnCO5yyNViwY26XJ6JDI2rl
wwTGB7ofJzjuhyrtu0g/ycZKh/rXSO1k9Gwy1cCMqxK90fSWgB/HEi9jRL2Z1R53
1a4Jp4hjt+ukNkqWL9N/vUOm9BTy8VR/F0ByILpulr1vp/Lnm2d6OWteZWUNtJoP
oh1K0PTDfxgrLOpWQIrI89sOAg5w+5JyaeT/dl+QFyx87SgGCkVkAfSeWRAbtcFg
9ei0Ox+xdpUAb3cmxYAqvq+JUkiVq9ot/YmtmzChYY1e6EPVTTP0sC3dyu3CDcZ2
qeBcWQvAQGL0XMfcdhqA4csjxpnqBFjekPUj/m+UKz5S/4ixEgRSI5iiRE9s8ztr
Xz3ggm7pV/JYtz3EPdurhi27EdWmQ6e6DgOIO39VvHv6K+lUMGpIRb9IuY5Qqf0w
VhXixAGjOZHEGcFurWXpGY2jKzuXEsrouvrUy7P3kotX1/V1XkVUFFcNl31UBQiP
f7h4rtvnfk0l6UvHm40CRuIbv59bGVXtTxkSuBaVoj1IgU9822Tt8QonHsoHJw/K
oaFh0+7J9kUYiHBraWbU6hn1XC8Mzz7y3IXcbDjJ95mTwB6YeOZGPoFOEKbO15PS
kNxA0YHnKtJnOXe1DfhSqwu1/I8ordZ5tHNpDjH6DqFVs7XmpOPR/kBi5wyZ2jwE
bYzPnIT1f/0XCIuosNsED7GbQqUkTzXsgn9Qs6oXcGeEPHuxRcSncHXtsKatqjEg
tUq6syjZrB0V4/GPCq1GCHsBATz7oIDmqTSi0nQyBZ1WD4kKy/Sd/IWcPmX1PUoz
wDOdNvmQtrfPNcOmvw6HHaHrNWSnLlu0a6QkRRDyoazdgnDQJfQ8CWjHs9xfbVWL
2PwhNsreuLKoJ7MiGwTCaepWDdGEDqHLPLn7vy0TEtkdyZjWScs3h7G4W7Mnkmd8
n4I8ZvWXr1cq4POmzCGZK5DSeSOqE4GDEyitu7Cod81kr4IVYPniE99XWrD/eWp8
2u/IK5jRjmGm+q3n6lGOF03mUi1ZrJi55huhYfYa4wd8HuFi0PxKjFwab7WAS0nF
6X81aA5/uPoqUCP/DAon5NIkvcP62g9zXuBpMaLUQJqykDgnRorud1difOIminuH
BDvHV7qbGtuEOjumBAj/DLa15p98cCaRQVejrLQkgpnzdfChUSYwlzPFrKzuXYj8
p5A3Er9xrYFXTNvp7uLGIMLQhb/9H3Hy5EoyfF11P73XEX+32nxq+sUXuHHNj8NW
dPMvAxQzOkDDSUZ0U4pp+zPK7JVt/JC9s6v+GkcfPXNTxOs83jJSJnxDvrCFqdtg
SpeZ1ZyaZ+pPwfYkQ1cGb0GOD6U02OOBSNYq5n+LBh4FL2q3kqFtt6D6WfgOHfdE
yXiJqC3e0ahdGcT7CMradvmUUx5TTUZ7rTUnQVA9bmiFdQ6rN5F1mmSWQ0p+gM3F
4CBoSqIWvNkuiHGTlV/wckzReRlzrBK84WV463OD7KCik10MP0mybRhSkz9wg3uQ
tW+8yhz8JyLDPz4s1xBCcSUWbhY1eFE6i34toqmyeVd1z6AZLnkPi/uJ8pbshsNm
uXEEn7uzEZVgXgpzEbQMy1AdAhf1RzVBJHxjLRZr6z86ubpXaofSqK1s6ywiheip
K/fQxj9FdGKYHRGv0X7/p9XFfMGlMu2KSam85sH9jBseuqRcec9sWiW/utAdUx+i
G4hT9Jh4na1ndT9ld0bwwYQxrwAfHGw1YPqkouRcyLzYT8MKqEO8/SLGWqeq15Mk
1SmGeHS1lKZtUPRvCxuQ/DHfoDq7IQhBVFrb+2KJr3vwNYw8LskhfI9lLH6V9x3b
ZyLA/+U8/zDVIio3lh2CiVpX9z+BkZNhD7kFJ2atCEGt/eOWc/jxOLe9iXrvObhJ
3RYpWfgvNuPqPz56h2tjzlTdcCN48QcDdNAyLd/gDp1dDv2o1qC/fRENkOu/ExO0
4OkbJVSA/5/ED8y5/FVuVX4HreZubPeA+ibfoItmkxvR11hRYYdB1/TJlmp5ZrRQ
v7uHx86hF6LRTWoHNPURhQc8aDJ4Psd06n9zopaQGxfEDNl1Xhm95ZBy7Q5kGfSs
sTzHDJrCKKy8ypC3VTcVIGsdsPZQX3hzNuObhGvdlcEbCxfv0AyPFotE1XikYfd3
oRjS81L2x9oWwI9hGs52pWpsZp6IMzlPtOWjME9syhseydQ4fPtk4LPk0ztz2/E1
G3tYD6Ts3To6TeE+006hM03EuR2XYm0Q/3jJdbW4wxq0gY4RgeHC5X+Y4yA23wh4
v7Nk+1oV0z56DRWjScwJeIFQ74mx/UPm2LuGkPqcVSJFRpB9tcyDSq9/HcjsADRg
+bWRrtDiZniN8NFyCdL5YeUgJYt3zL2iUxvA2RV6UqVP4RrGllh3SIlO08wUq8Ef
5PiG/1IJPFDM2TnY0o1xLe9E2DqKjqiPoIK7n2Xo6Xli+Sh8YdxZWYZZxP/5IIFK
W55n5Y2Fghfh+99PAFHRIdcM8o2Df6pIq1xP7WMt25faWc8ZCAdIXv5yoDqEKkrX
+iLjUCglOLR2NgyJNcarqK0P660bthQdeCbMeZA1aQQ8TLpf7ctLcWus524FLkDB
QXX6fCeQOmO9kfRYLjBRzjNg0nhfu2w8bbiPBWbzIbHm3b/1rqqQdY+gvvl85Pxd
ctDID65hebhOn0DCBnYf5zc76o3qW5CBopEwqEbGWnmI/GwtqVf6o0IQiVS/e1Ac
HljTOn/aTTCdWYgfEl+uAtyrs88wLbgWt5MbrBWROcfGKg8+RMECvmWAKQgnjLrh
684VgdNSIJ22gytKwPQOKx7Tuc3zo/FYIHi/t6a1OnKq9AhhuQ6fyIFFxmrxfwdM
BU2x2T0x2UNeh9HIA/6RA5svosILF4l21zRPbjY8qHmufrj2R4qX+HIBeeH//OD8
KGpratllwI8oojjuKhxVItqU/278yt+ELbONlDfqI3n8Vgvdh9uBVktjVYZQwHLW
YtoqRyyEmwogw1hRtHVYSyY8ZymOrtpz88/2khKcQbEwV7grNds5hqXEwspvv8uR
9MXcCPmb5oyBMkx0QLzMgzzayKjhyWlXry3uMvvo11pDd9Z2NWskkKrKTYH98oZ2
zjvoerlwPuhPa49F1iWxxFFCWqpVYic4FKI1cIRgOrFuIQz0rC+NxAilHVfonypy
/mhXbPe/MCdcQvqpKlfbqvFgbd9t/85Buv3gbmXe8/ModuZajb9PC+g1cZBUzaRf
jMpExyp0+DqyTLZ/t9KAaHr+S0DoRFgmvh8ylvcbQuqZpk51+Zlp8MaCQ25hyTyU
8Ektig+ofz1mHxYGtNyEDCxBM6moZPnstwEnOtKU8bH2i19KU5oumMW5tDzgy0sm
7YP5z65wGrb8mZ/zEFqLYjgpyx8CDEN1+UllT2V0OU/cUzcX8yHZ10dfIJOLQjyG
HlUAw14i5vGab0hoQWOG/MQELgpTh7bkbykFk1B5R4nlR1FcBJ4aEjel39Qy0ao4
i0nDHfShBsREtNfdy5ghxzy585ruwfTqrH31XEUMVDJB9S4p+7Z2izyk7WfU7APQ
UWyeb0h0N8sH+1DnsICEEJvgzjv6MHNoXOry1CAlVfIxrL/b4w3wmk0fMx4dptc1
5/HB7YdFw5r7CuZ3UkqHMp+4KEf5qp3He/AKSIErT8UsmdnanvoIpXEVIVPX0ebv
P7iaT+UV53XlSrXUGE5+iqqvg/u0Y/UH1H+7HQyrTcIezWDo2RxIgP8Q2bruzAve
aNkW24ugRg9ErlzDJV1ZqgbjD4NKWssogDk91qE82Pj0h62a7lgqKkz1YyV7ZOAl
X2rdb/q/s8hxIvyfLpkJc2YJvL0QcTIi8O1Nldb0PQM/4v7F2luHknx6bDQtBfbO
G9nxtokxaeu4BjvIJXXRbHT8oIuZ7c8d+th7xvOXnAxSSdyhF1zGqeghurA/Ln5k
AqXCPJWIivDGrbw7lwJIgClZOyotd9Eg0TrWSpVgrwp007P10e92oUPMgsLb5QtD
W63FE9RY+rkwhNmIUFeFJPPhne7TPz8Tk86lE/Qbkwnm+hPZQYd+tApzWtA2BpvX
IiSAAD6fimzpxCQvX5gV8aV2+iS++NpOp0YUYIpHZFWHwrdNWdLBA3x7IuvriDe+
/PepRy/IFqgCSdIwmAuNgF9Bcy8es8ZeUWgpSanmCFev/ytWjCZHG+vUIa6xH+BN
WYvunFVQuoSaGY9EZqq1L1lADyY7+Wc79/bFHV8XcZXAGOSXVPs8YpGsOfwLMUBT
6WL/Exl+2K1JKUGzA7ubPzUs/GrPxJmORm8+i70KlCBnhm+S/zYkPoaribLC891h
TfXaYU6V+K2amrZOWqh8HFFf0A5mydtZrvGm7wJ4i/cRmAw/fL8NuO3dP7D5OGYH
fjTtQlLQZmHcz9s0Ga30uUz21q5ic1ymWKXDXLLb8fthyCI0lQxEiAZa0YrgLVpi
oym9KMZ2oyhAbgSMr4+gvTKiBiOvdYlLflv+OgGne+m1CtXsCgcBeQKy8Hvm2533
adsJbd0maDRzyP/In4i8HiOEp4om1ru4Ph378W+SYFwTXI48ZwKMwFC31cMvUwi2
k8B8TW55Z0AVAb8fcX3c2+ypD9mMQkxKgqg6c7ct/ijuoFxAsZcpE1Z28TU3d/L4
3IYn33GSUwSimoWeg6zecXEorOGu1TTj0zI58YoH5qrLIMKmDXf8W+jk+RDH0QK0
65fS039u0va7G6NcB+eOBwOxlrKPnbdUjTD4gMR43xE6L/K1r2OsaPFFoL9bWSe2
nz/DasVpdLwYLl86r+0AcbmrIbV+wteEvkJPIzSosw9ZR+EEDWZMpW+MNKxKktE2
SRrQ8hoW6KorQPehk9wonh61/6XErTiF+2Cc+4n2RCm5Am/DU7n3+KHWlJ37J0wU
t8ZeSGSKR/45cn3BTxpoLb+xpINCmm1gfJ96Y9/3+0S52frhXVizV60cj+A3+6bl
RPr+1Vm2AGjvrXEaT4f20jVC/OF/qqtk4YEPHiFs6KHm+RBUHXfrCLpAF2vNoA5q
cWEm6Dc8zOOaVPQQR3h+/XKx/6CEE4eDHOk5pE6dg+jwpz6hhaRIV5uMq0/LgtX+
9vl2OZGhYb+Ce801dMNNHBY/ldd8hlp94YHtMeU/LCySv4TuX8R+2pWCaZShZxrV
jMXujLbkrx5aFuFrZflsqbhmieCA11RW4jfy4WmlRwXcsQAWBdOyrun+gK1RJRG+
Fybj0EMZqYR9m27Ubx9/jXY1SJKm3Ap6IekHbbBg0QkBN8836Hz66TIiNFj7Z32J
ZjQKq33rxEFahmzEo/oGtFSzj6wqK/DonaZ+4k5zR3Ies2XSPkvLVqzouCJOcVCz
xrVVLWokTzkKLPobjnm62IRFPrZAkq4N2tjJ+L55vLoJ7pxlJlQPIW38tQMG3iiZ
B3/V25dZBiXk3cfIg0iQJVg4ahe0bCw1bNtpwVM/KK1fo335EvLgag59S2dPp+HO
XouI2C1HMJLexEzCJWbDMMpgGIYGFCU5adYypfuF5zi7AjmPY7EXMyrPnZaSuZl5
5Sbw4hGOHBxQVXMEWp+Y0HpPd7uCpY56PUgzWmnANoR+5yI17XQyxHiA7rXTrKEX
YsRZf47iGbVD1HKuY/Ux3/RLDVtaSItDOMowD3QYHp5Hk852K1Hnga/1cc+fSPl7
vpafKKoQdwtOis8FiSi/2r6aMZPbBzSrRVPbx3PlOLN/ponDnSUXFDcLxE+FnpJ2
Wq6Y6JukK0PZozOHZYwQmShWU+v7pkpPtafFBFgiwXSzhbZbXvjJY05STneSs9u8
YlItfVv5SjmnCHe5nRxBIQ++wTJtex9yrTgTfTdI3bqHZMFcdenvldBjrC0hPpIT
x3pvt701vX0xOubQwkKUQNWtMJsHk6p+lt0X3S5KfvDNoFv3NzpD8snn+ZUcKvI8
pxz358lNEcySciFdIu1TBlqFFuKU2+nFnQSW8AS+3MJIo5Z4HL+kuTqWFKlxMGCp
8PszCP4MXOxdIdjBjBXP/DV/gZSOXCZ/+RPEmRFXKFKBuLOEuswfu77LbMq635t5
HIaCdj4+d5pS2Vqjno/bP9d3Bj9Oa5FU5o9gEa4zNJZ7Qh8w1K9PdIhjywtuRNgp
m2GZw+RaAn2V+Qnwpa4ux6XRwRip+PExEoDQQ4WeVdujI6fSGeSh6qilU/H4cG1I
k7e0uwv7bURNrhvD+x744sp+PIfjh2vYrJlxWSJ13nV9R7al40AD6F7FulP8IAS/
h8/tq+vNAeh6slszolom3Qd1m6khCxvlVTzslzyFDaZsjlt5coTa9PBZyKlggZ3N
qIUPKu0hWgyFc83SEhdtkgAgrbv8pMeaGyz64nYcBWS5mQiwV1jO6yp8IG9o3Fkg
1epmiTLe5xW09fbvqhkbw4SuVM1xlVywkG8YMVd4RY9BvIcf+zXE0PthwXgJFcqd
OBQzcJCSivYmaF5RKIhMJg1Qx/3z+vnM8OMeHyUgHuAASmbT/P6kw3WIBpKCzHQH
mjIfnRZeBAn3URYa7xjAHAbPJ4VVfW+Mg7OezHCO90Cp9lGWL95gkyBPwPGsBk97
hz77gnnpdaajopCQ0UwwRA3xEDzs3RZg7q669We7FlELWf9lgXMiGNPdOfxyZ4LI
BUQfp+QFblrr0zWMYbx//yy8R0Jf4dzTMxuIhsYSkl3zTj9deoVv2ARhRYblIEC6
aQu8ojoOcJG3WXGM9on+609zO9Lk1lRKYoqBu8PIvUfrK1oOZNGvoVrzNwdvtPiv
CbS7wktUhk7UqS0NpfWlfHRD9epUhbOhoAHn6UnSWssaK6yoSyNM4k8vojwlWcxj
GfUamI1Ujp8zgSPZOjpsBIoeloDNYVlVUVU9PegnkQ/Cj8GZg+bdFt4SMdYY02kS
ost5BFeF9YWGVfgupAISTMF/9tNvCmXb1dNGLbv6AId+xOlKzv/21cZXpui/EizM
ifj6uvqmoxToaHY9avrRs99yumOfFQDbdlmCdK/s7VhpabupmQI5Mpt8bx6efAHg
cZjsjv18Aj58Kbn+XhYfdf2C0hUbaYSq26hILJiQ4OqoqBnJRahFcjiwgu8n6Vh8
8EBqQ5VuOG7om2SFUnOIpfh+y8zA+HcVXMWuNAWczaB+QuzU9mUM9zvKLsoR81kK
rpKiAquKhvH0ra9kICKny2qBGqhXXqvFH6clO+38BGn3GY/CTj8Oh3K77ZPbuIHc
jkqLEujvguIQXwc20tSwT6pVKEf6ZhTSaVXKqYduwHLSZ0r+OuWcPUde0bgl2ND0
W6W+/ZKNUzZLADzvgJzmxjzLP7ioUfsmsGh65JsN8YMKrhVMUzrUAyDUeYkvw7ij
64SKj1MZy0Xmx4st/2t3MRlBI6RVlO8pdPOJHgszY/KjW7Pa609szgQqMgj9nWYn
Eml6t2EXDze/49u62lJKA20MpeXVCSHdb5ICB8kRLQH0OS47+lRd2TtjeAA1YBwo
`pragma protect end_protected
