// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:28 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TQqiNTVujn4ZoX9bNDio6uhJFVxggL1klG2RU55E7XHXvaNNGseMy9mecZ7IXEHt
9+/WsYFtpiw+IRQyWLl4BoFRaMuDJJCiV8juP12vJboZSGmaG1Prp9hLear+d4Zb
OU9zMtOkK7Qpt6gx7S2w2sedJuxddSNOCq6v8ItubQo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
BHWJmh4LnB6ivnknH4XqUcEbFXNV/PPK4J84ManyYq/q7bytyw8H4V7flWhoCuMp
vYDtjLLV8vNPNauFMa3AJdU7Z55PhmCJztkrttkqrfDvyzNcdhuM+hUImpBiLIqD
P7p3RRyTMYIAO9gnVtxZe6VQfh4FjiHil/RDJC+V0Kl91hvua9R4hGwefVw/5ASi
YbpfTmr++bMj3NgBug1Uu53vzobcA/bePm4mn7G9cci49dgamAFjCyF7AoMnkSg0
Mz83f4wWCaqIL3WPvur7KyL7ReFFFVzkJfXzScqFjJwUdAzZkEFU+No9LRY9HL7k
tOd5szof56UsDBkB7xxPDo6u2oacJpOugczRqd0viQNpt3CzuHTBMbwugZjfHzEG
wdXKeuBpPHv2a+gOHxRNnH9xPIatyNyn5yUSnsWQ1qCIIuE78GtcmXtQ4aiMWbZ2
xC3EpZcjzlDS4PBMPWma0lxFr5BY0E3olT5+TojFkZ2jm6KFPc+SsL+zF/k69NZN
UGFmQIqyXj8sUSvf6DxEs/4z9KSpflDDDvb0d/MdPCyf9NRRI8iTpPoDeqN9ZLVv
7Bg4TVS/SwSIRCORdxv80l6cq3K5wIA47GH+zmhxWNFRnNC9Yuy0v4KfT8Fcj0yP
LYuDuj903lmop4QSNQh2kKIMmsqKKjcPetiYQ7IcYBKQCDFwQCPJrcmzEWFArsLJ
cRtJKul7B0Weix5UjvIBa1xv9TfiTVKAEG644hZEFZMRAp+uOEmgU/Iiizw6liOb
XQPPyMTVKXFJ5Dh2GRELRH4ECHiO1cIlGylP5rPkhU1HfOLOLMkSU0G5j+FJmyZY
/YW17eghDC1XcKSAEYiZ2d7wEOmBOPbzs612J4bz9UoUtcjVMVHm3kklOrMlTjM7
s52/fYUG5CRqVyo0jwNLDOax5qMDwepgYgRSgCYBkrEocAtLpIPp5uPJzs4Mpcal
/n4TKpbeVzfZtgjBwm67k3XsJdQp3KOcVPreCAv60fjSCHzvSoEX3kznvbSGLTGE
V7Rh72Sfzy0XUuueUx08rYPHj/jfNmAZq9fnvjUUX4MAwTHoT1uKDslBc+/8R4XE
JLEH97WzuEdOvYGVUMrD9JbehKf9SBlKuHj2jGa0UNSvQCIgblZ8PxZBl81mPdgg
Hsf4es9tT7/oRZOaMmnfjelhPEgcMYpSH6UEJXZDo+EQTSSPw/3zn5UmHNFU0V1n
ASGbMz5gxWYWo7fgcO8MntmGYi6tYutZf7V+rFgXvPpAoBxZB+6mu8Kqe2Ht6z3z
7gofcoej6r3eUFmuHMdP4ubOgWjkh9xBaWCq4dukphn9V4QrPbIuF8Ww2NHHTcLe
WUGVUNuwjR0pzmJH478wASWsAjsMXcaLymEvcO2JhaW1frlRt8YuNUtwsryQBIfK
uJspCpTA3pMTqjMXjxzCe3+zkg1qBijTrinyCdaqcezH+soIUByx54wFnK4bsdHP
0zzxmZIUIM+EJrTdMzbzFZPwzDVveATnXMMRsLXRVxJrEJdxJFIVfhjpvT0QQA3n
8h6m2CPkSUWMYo8O9IUmmqGJ9aQowluFfq6W4pQaPUsUBYNhOweQSyh/6jaf6mKQ
Yc1M6CNMin6LC2PG/xf2pScoRQRxBaZ4TPbmfwPuYAP7YOYPHy0k7gFGovvLIWqY
KLz0VJs9XopwNgB6tke+WEp3/jwWhEutJh5kkECbwwG7flWVWWu5LSoE73Y05Kci
0/9dpNWdZy0h93lzbixUQrowzrT4bfbw0YoMYKbU+9v8ZCeKN7QdZAHnswC5qq1n
z7Kn3MBA4bszjK+SPH4CetUObrEWix2XaZqHn/KABVBDlJ+Q/5YwmlS+wdaepsYr
+eJDTKd8xRfDqlkhXJpvKqPKkCLYewuk1gg4jIpVK5djRVKlcm6/OeLbM1Xbx9Ox
7PKf2IcjGyBgvg38HS3oPz+SO65n8xyHLDdmlUj4GvPuEfjxxgXNWv4Lq5Vh5kdY
O9Cd2Wq9/57hM1yZtwSaUrMOPHMqdrrbUig19i8+k9SY0daRpjq/++0TNS2BG7nf
YHMbBXBNp1qQOMjxwEqjs8BfRCGxb2mQenCzTS676w/hgaBBu4bTeerIbzsbLl8A
Z2P0fKNohfseNJemLrg4v3M6/UasaopU0+vaFfMSuRi4WhqJSjrOjydvkbClkgbx
VVHrUwbchABbiBWv0KReJG0bFKsLWABKAXnhJIzt3vsgW6gjZ0T2sCpJak5AZwG7
3ZV630YVS51DERsoabd+OT3MsYGtvN98uq8D2RwZEQYbKo+6G5vx5JnwrkWWlr07
4X8QEyHRumAxjCTY5SFKjg83KY8RUvNxnPzDX69ciXi3p5UCetVbwpN2ACwfD+q9
gkCh62Hm2RnP8wuRdfNEyCDhmYLK3tsvnF0OmHWt0z8IDGJPOIb7wcuZ5ixLC2Io
cUPtUcODVMBxJGlMggq3Nt2gRoTVXjP5ckOgC5nBSF/EhjmeZlXgMqWkfW7xHSeh
a+W75JAiEU9j2Ewpc7a1Ao3R7+cpz+Ej9OXypLfpMKlmKZXVjxq83EMaVShpM9uz
M6ZKbvLWqg6iX7EWGqnujBjVwvgNTEU0FxZ646Y/CdQkLITwW+mI2ThzMrb0LU9e
Ish3zOdSFyPADKEirkZBcC1HL4aIrYdF3VD+sCGr06Qv77Xj4Xzbqqy4FBl+vglC
S8mE6MhAZM2lJYl1xA98+hDccBS3idWkG6lgoIfQcLSnTTemr7wccDU+jD6DEKdw
z1dAGowg9vtfJ1RHiftPTwQ45Kejpzj/K1aVum7ml/Vrlx0LWzPBOOe5ypbC3IWZ
vCtqZH0pUYP03N1Vfe3cJRdEDcBsqYSf4JCCB9jtmwxkUMfeP2qbcXWnlWBSs0TV
cvW4M7RJDBGhYaX38bD8DJNoNe5Tzmn1hk778Yue5FPP7NZZYN8BT4K16KxLqv/D
zHrmNUmdAbEAp6W5PgMoTDzZ+3t3IaE4y6DTggIGapFPbGGexCkjxW1jKIASIGiF
oY5rpWyfBxo1b2Ezy28w67V7X8/DPM3P54vykzabshF+20otmxaxN1Bdq36S6uaw
EatjWouowbrRD+lRHx48BQjuHpSS8jdqm0+x/K53ZHjCIZKjQ1mpYnv9o0jIts04
63yZyOif7geIdIeHy1Ex16v76y2TfSDWlyWo+r3OKsaR9NHrX+nXHDVT788A8xfB
0C3PBuldxFs2Bdrx11qAPfeoh8o9a+3nxNaOBJ/pxIKEgagLk0wyISs9arpfYM/7
0oqcctywa9fu1ngs+RUmi77/LGmYES37yKO/Qefspn2R0GQ8qsmvFS1S/1/qOBI8
TzajCcabSTDslpxpUDRHXu2Vhl+yvfUFXUeeKmtT6TLeGU0aIENWwKs7uX+UvrOc
RLG3qpv4Fi82qa+XoYT550oq0xx6QrlIZwxZ3u71losPDR0Q775uq3QhtDBxbv/F
rkj7MEKcFdztlkzr+6OrHMmOPGMhjzeiSIkzmF9GHC/96vrfxZ4/qk9w1CYt0oxf
OCLW1FqOLlf54780FYJCftP8QyjsV5ATcrlPNURT+MB6JeoyxvDNUEW9aySNyv13
4MUb0UV4ASGe/I6+z2uKGCVvXeihoM3U5Fg/ejniMWKXXH/C1CLoE74OM5t0VK2P
XKvDD7sm69OckNjO6QtO2kC3R38tPDxNjfaRsIc0btkWZ5JDvKYfl7UuLSwEFryT
6HmOwqbXldb5IvUPMhXUXPVd7Drm6vcoLxZW79l//Jq39UYUCbN9QRRnwi6PiQni
oEILNvpQaWlU++SsWo6OEAzMZ5KRR4YhQdyfLOLZciMFDmDmdgsOEV3M/myNLfCH
lw1e+Ag0YaV/i1Xel3YDGNbn93crlxQwfL6ysy0YBZzRQEIEXq/LIz+OhVnAeVMF
skyemQVP6XNwNA8lhAeZbl4rYP7qkCv5NCG5ZYLoD6E1nUOR+NGeAAbIYXg3PtMZ
v8Q7KJYuVuP0kaewpDc8AY/SDp8xHgpAWfl/aKI4WWVfwwx2JKpVHBCKlJQ9crgC
7BjKEsAEEm5T7rYRJcp6WQC626CruyzZbuk3TEgrrOOQl0KMXeVAPFQaAEajLvLp
dtipl9bMaQ5YdMaiSVXTjoKIeQaqOfWKaOLl3VhCmdG0cXlFbRYkaFCPtUDeCQwG
l2qy4YFoX+KOe3Gpq8+6UCy/1UdV74z1QDh9Sp4OpU0CUKG3oNA2PM43hVlfUOiw
dZTerjcsPB1HX/z237/WXkq0SJHS2v1YgDiE/4M7sflghUPsxIVVQfUHBSaKBMbF
WI+JoFWDSCbcF46aspRz3sdB7s9HdtRP5cgtgOKXdIDGcZLjyTtymMhid6nYbDPI
ottjPJNL3Vxh888bAIp1Njrl8UXRWWT03sAilMOQsronIB6bTRXClpjDglJ2U7rL
PmvJU5CtZxp1yu4FrgkVQaGCUr/oNth5dJLt1BXtOdvkDmJxE7McodZbnihLRMI0
NtB2iGv25AqcnqehUJBDeUAKiNCZuDF49F92q2FMzNWmLvUHBv7tMhdi51Dn++oD
GP9+F8A6pDDnUsOLpJ+jjbTFsp84LsERqKeYaNFatSXrFZtzf9WNahHnBpovX88Q
oTLg5lYUNmOYNbFQqK6HgVmagsLwgIYek3PhBtvCT0/3Z0rHetfhxT8KapeDzOyA
jCAA90Jpl9ag+2QqyGLxuhTNlrTomwN3jS3R00AW1L1JG3Af6xuWWCItd7O8zVQl
yTZVFZqIAJlC324x89+CGEN+b7EVm8WNiCK2OLSMK2A3i9Xx1FFSrb3HFNTJpV+l
6gf6lJH+z+rbv8HXTICQegzvZ5FhIEY+rax2Dsi/FL6+abrjqKdA4uFCGbeMzKKk
LRnoim0Oa+JNpcElqe9AN+tUS9anbiHvrKzR250+nV9YRF0sOniH2XORODQkkdkt
JkmJ5AOiMsggShniqp4Z2MwQpnug0cblmdtBBbVNWfa2IoZUx+RkzdkIDbB7HcQ3
FjXiLsJObUvbxHl8fVdFbMKLMMhVTpLy76B1/22SHUarPWCWEJ6Y0OQrp3UAyl5u
7d0hSiom3dkBX+1/G/xjI5pqbm12apGQ1Z9fC76YrH5gvCXqKveQaPocfzf7P6PA
MB6/5QDi2P4oOuC8RfyjgdBxVndZts4OSRcf3LUt0lGt3GUGjvVINy0K0FALbRsU
oj6XdM8jlrwR+PcUyDgzRdEh+6ngPiY3jWrCv8FK2g7iR6wXnpHvUXUPJkXkROn3
TVXBuE5lE26+4kNkVzwib+Z8qWqxS6Qtwabzmbp8QDNu07/a9gro0rkdGPjVY0lU
B2Zp9aJIqkcd9JMBq9t5EbY9/0mpnZQUAJmV5dRDv977CjcetTGiDtgT0enT7gJ7
f4LUwqhPYnIuxyKW2EdjVxdWpUrN9XSErZGqirSEiUUl6JStoHEkmwseyQS8OBS2
BP6vHIe/hi4IQpAMxD68uuxc/KoSUS026w6F/AB+2CbI6kbDwmavygPW1Xl48QQa
GrFSjiBP5bh0yJzQ3CzPlyOE3IL8MhCbwkCWYTe0kV6uN6DbdRIo9xqC1RSA8Qcc
7rFr7ew3kmkQ62a6wOv7Oq3QBKqNeOlx7RLF7nC39WYqsY/SdBH+VhEZywD8GrA1
46m/ng/Ld4Qy66vj2FOmKxanXfGwMXN+yai7KFykfYLzYbaUb3QrHZEFnYM2UM7x
lOecswHBBYt+F5mE7uUP5c+JRdBEte9o/boV3seICoiy42pzNAMXYzPAHz8jyLwE
JyX6gNU/1DJmzDD9suPSxIc9S2G4c0pw0j/b6VP+SgFtherXqED3L1fTeFoz6JVL
/ddSRS5ifFNnSaNr8MJgjDbzGzMQ5Kk3yYanAlwQC2IbhO7b6RiMNem4+yzbJ75d
3TtiS5SgieixkUqBBHYpUFd2UnR/nRIiffdWM2drlY+1hI0QoNh7NDsdmpSqN6xX
Vi7reQwNtMRfGwSAb3bMgOW63qj7sJYg+Z1T3QMLO2YqYAtK0dWFFZK+ulALIdKQ
yd7UOIrIZAkMsRatj2rCv5cYg5/LH4cdjtc8XnjNocKFQdmLDXa+CixgyOHytEqg
fBqz1LioLJQGf+j7vojX2C0VCfin46TGjVhj3WjNAy7DZ+H630c/MWHryE/r5Svp
dzzx6HxS3ZwTDxL6w5W6vIjOsOFs6UxREzjPx4SngsYSZpDIKwPIk71nSFTIg0aI
DQa9YsY28Vk3ulOD7T+XJrS/7wIavM2Y3YidsRUY3NAPDUiAM3FQxMKPPtZPef78
6Xs+TxSUyGbvbaqWe0LIR1yt0MrL/uW56mCSx/NxsKFrevF/YFUDiTovX6IS6D+g
aZg2G2z/mEDCpzZwcDrFrO65CXWnaPpgB3FwyIGnycui2rwqNDyfYlmzYeMGEHRl
5UeG6Luwmte1hRjSI3ZBSt9BhLn7PglylEBzXg4GKwGYRbN8xH2f/e9icxs5xIw1
rGjgk9e+/KLOnICISTeyVsaSnjOu+hY0uu06K/1t1F0GDzer+7MEe303vCDiR8qt
515jYcPk0KczE2cf7qtGkTy808tmQQkvlzTGvXN26vrYNu6jZiyrakccTAsd2SZr
BKYn2dKfPovzuEL8s238872oR8N3DFXsy6381wCpvMAdnyJhoQ4WP1hpUPZrEVBe
8zFcjF4znw9BQv2vOwAGrih/boaxAp6GCig2XtxuskOuiFsq6mEmu/KikscNrdks
GDjcsAuKQ66n9YcCBXI4L2Ty7rpRv12weWuDeN8nwxnFvUHJD2dXQ760cP5lsBDb
hbtZkCiG+UEY6DrzLq3c/AEmGQ/MqYdxzYbffkl8GIaXWp72qBEB5CZuzOCHbyEB
A98nuLYfhi3uQmGNEgwW8UwYwzyfRm+xtssAsszkdt8V+QsKqV3ipaX6CObjwyty
snBtWs9WiPvZT29yxLJV6E0dOeh98niSlCzIV5+yrAKX9Uf9J3hklq9t91WB1hRd
12MYPu1RmCSeVYHdvAhCJpTRe1dlVI9PtWJKLTZWyWXV9viu3kvUm3g20smD+mGY
pFJqqtr3pzFf/ebJkH1s5ZJEM4WsiNS6ICPogiGlGfPSXUUyy4Y/QNUiBE0/XHHW
5Kc5gncAhmoUoMzctwTbiIU17fhteK5cSVCnksRk/jGmX+6LyifIq52ANpMaX+KW
JSYUSU6ETKOiUQenGioAF3v+1LK4Xt/F3g918JEvN5nWkCUVz3BQUkx14vqA7Bs1
Uwb8HCexqMcE+WJJ3corjOCbJAHIFwMy+nPnmlrlNJtfI/UAANSNkzH+YI02LTHQ
xZHKpy5M7E05wyNwWirOGJZES6Ce8GHlXFv6ItFw331g+QXAu+KC2T4V+ADONmKT
x7wqtdHwHpFcbN7qoEa5aBybVRf4P9nzDjTuK0pt4dAiWoMNhRiWLHqWDEn6LCsH
6rpUmzeRjxv6O5G5j7ddxKML1j44nzgSeYnMvVr8xs+2riA0uVIMKtgKe7Fs7+gm
IJDLEiySvnwlO7EPFH0n/AeKZJMuAnd+nchzd/hS2PpEvauOqCfLZqTanBBvOHTq
qv6d40h6P7NCaLQ7r1dscuNCNCwaTL92YCcDKRPLStO2gtkI1v5O896wa8h48HDB
w7Krh+A4QpOFiu4qvY8HOEkcU0Xe0ei904VcbZqevB/OUORR+/J3hR0JaWA3DkkM
iL92F/zdhFMMVqxiscRbyohslCqbuVEJMu4O8sytVjPEMLi+jfB0n6Ugk96rsX2e
2q6fJ4pVMcV+H/XcbUlEsjr/xTLXmf9dm9mREby+qXV2WtVsZPp+1U1ro7a9BPN7
MrTHsea2+h57MxwBhN5aQjV2fMnM96Kv545m2g4SpFvhxlCU2+gx1K5QyVyBvcaa
RtLybT1eFOYuyjt2Rhp5rz/EjM1Yk+dkCv7LhvaVDRc4WzcKQRtJdN5bUChUarGJ
xnzUK7YwA3lYCeZPTFHBJ/xMKMb30hX+DQFqDPCw6TGdE9mmEMee4Fp3IbDOt250
+9Twdb/FqqEeOYLp8v2N3ywAHWFc3dqSc0gjvuNqzgp25cn3n+B7+tnhTDH2U7Av
xljkNh+pkpe47jSaFrSoHECEjANAhhwAF+u2ZZ45tEJ2McNCXDqaaWerw7OHtZfe
e6zppZmwyi/8BZJxeMyT85VkfwET6x5pQCQt2WiM3r148ENlcLp1POYaAYa5XKmw
aJX4bbgh4FcRSG9BZE86PMSE0jyn62HSwo5iCLQrMtgoDbExYihL3Wl4iJnBKRhA
xyh82i3ls/2YZcvLKlOVTkErsCCrlXrbWDFa/UsoVXCSgcmUptJxJCirvopRu7qC
maqTGmKJ/sg+L4+zRI4cQoWJvKafrDjqqa2Ca/7awFwgv5/yQNtGXjIFf6fmDCxt
Er1lWzLI90+YcQMjJQKbYz0rzfgw2Y90cXbxsK1KsRnVKaCMt+tzO9J+dOFsTRsN
AvRWWrD7myRdMMBZhLVuRp7slkuY2kQ2u1kkpjzUQfU7wHorgZwxLjb3no/28Lxy
4LfJsbISM7q34cOS+m6OgdrA0ZC4BiSMgnNB5v6kRRZdrb1TpI2tNSW64MVVqpp4
vRJWmnrSgMFGeri8PmUb8aLxGnP2Zz/h/gp4wyACD90WnwWttvX8WJnM34AiagpO
awVKhcZ4u6aAjzejd3bmerz6GQ2qNI04pbGQF22W1nVsVUsRsARtYyr+KiI2arGE
pmYN4udNqgB93NTnIwk1wZJtcYP26YvRGKJtmpe+O8cqYR6/5Lc6WOlwbAQDxjPd
tj6di+fxktSjA4kcs82/zS16vD4oYwnXF01gMM6X6U7sIQo87JeTg+f3XwDh54Rp
poPyPx6PrCxVaswKrIrWeipaWPD8TPHsEsuxZwZQYYcU5a4qruuvKrIpym/l2YrU
Q9oBJ/NVCrdh8ieIivZU1BmUjY/5GU2cao/IbvJWHEZd7t9GVI+5pxFLNvdRYyZm
JqaOZRvQC2RoZOuGnizUbGK0dPa+VH6a9V9gtCBFs76pkj+4cHYsAkyD7tjON0WB
p612FTMcIDrVRuzIRqu8MmpDfjPKrz9jTWNDYL8IfG5dADzJ9v9Y00PR8JReqbZm
RlG7Wgk1cvAd4avNK8s07IhHHNu9MECuxBSod6xVtl6g7i3uyGnZm8zTt3OAbIrf
wDvyB4cXpSU55zXPFnV9fpKiqVEEsdF0IdplGB68hpTDrezRlKR4h45SCzuidQH0
bQ4sd1fpxMTMsdgViMKNDqWR49f+2P/yrMbB57NK4touNSQEb9Gbnw+DFeCwEbwN
9lZqCQa8qXBW3sApT3FHDtxVH01Bq8gvg3mGacMH8y3Ooh4f+45fNji9U67ScXNX
3rolq6hP7+lQI1ZQa8YVRAxVUANRgKUuQPLpA7ZmHWwfk4YwGNyRIJ4Gv8JL0ASr
DbqNU8TeIvqkO1EWP58IHK/Un3cIOO3GgUXhCq2CME85Fth761+JZgifFee/PS4Y
nI9JrxwME3LuHtWhWbR6gl2ml8SZUzC4mQwwZMQYzMWOwysv4dRSVmdnR2EO8Tpk
jHghMPdwiUFdoUfUnnaeFroKRigGgXJkCGVRcjWnpwFeD1vPZWvkZPXCO00ycYTu
ouHpkv/A4QY1M8K8+Ccohz+rhRrC0uD047oZOvS6jzcT49v8ijIeW6d34KXXRKdM
GveLYs6ZYEZluzBatlxw2U7Qj6vpGbal0jLDbdqo1CvNKJG2CLaejGkFFcOWPZMp
+ZSewGPXCuLdEgrn2N+YbPkfOrlERc+AV009mz86y7V2AcWHp/9c5iV9eXq9nk5o
zOiTbIbjuozg+bDaRgVj4lKs1qMfevVlmUtIr4ERpyND96UZnd4j3E14TXSP5jpD
p5pb2H1gZOrhL1XwAL6ekSxuw7Lop+DDIQUK7/fe/alXyxH4L6oOnvZD1LhmyMLe
L8mw7CLC7JKPl+/WRSZ+s03S/+aAo3vXSHHLehYLHVoASQF72udmYjcQuwrkLa90
sPqT/rT3/yOjnRLxpcLtLaAoZYo7N8PZkXRo3BFCVqxQdifzSQIWCo3Ci5b6Y0iD
WMdC01m0WiZY0mR/g6HrR3M2m8IPKwM1+rCwJtZvk7MXXF/BOzNZXOSYXtfAsP68
1YYhKlp/J8VdyLqPFIujCvHI8p462scCRrpD1zq29TLkcwnAYehNATBbOLDDVxCk
R0RceIapFSTQ9Ax6ylr6f0kQJnejv7ShvWDpHcETMD1A4uq4iJ113bDAkfy9i4S0
ICWkmaCzNhy0y7cBN6mUoPQschpEl6HCysiyOdKMjCcDNeR6b+a6URaehLIZbBDs
yDCWCAUO00NKF6nkakeSjhR5/vFLehqVWqFpJITSQZgIKnGmBIQZOB8sX6BMB7cb
3VNetNDzjKL3LUOWbVOw//SI4Vfz9uGWjI2NmYqOjrvF4vz7Y1OR5pH7qIOE5iSC
thmDu8jqd94NqBeMQDiYeNJvaANgv/kG0Ihj1ftWLp8LjB81/C+4GmrQ20Dt4ZGL
zgfA5HQPEFJJgtCDyQ/VcDTs4kNXqdg/f5yXSc+lPfZF+/nM6k/KcMY51dR+Vctx
`pragma protect end_protected
