// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:17 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JjqcII9nFr4kDM0oMJfTe2uchG+Xt8cVPaGHNcfwmy+Xisrp4D2ARnYFh1uf1KB7
fiVr/ZxPGHREdhmLjz2p1l6fFllfBmCrA7NC1Hn4zBajlqLPQe7R/ItFtWf+QhcI
fZpUOTevJpsC9FgFzqotY2rx4QPAihMTfIe+DEI9Yng=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
SUyia7zLc3foEgrhkkcPfd4O0OZBkHVAQMdDtIUH9+nYQ/8bMdKxGA+Ws/DkwLAe
vusaw7E5DI2f63eH1hQ07/kSPRJVpietR4T9RSrI6jF0CBJdeEeCN2VHdz/cN+OM
dkMcaB0rk1/zO5KBmUxgTTLbpniAvQ1Av3IfRj6k9TL4V4gtqYAqZWhA9ow4+bl6
6X4AETSyDz6A+K+z4rI5WGaGN90H2Wu7GMeN9RmnMoRnaGc9wX7VXvgTigCORF9w
bOP4697RkOgcR/gmITuwYdkMH1k5c/cvvsKuRovaTUVr5kv1oS2S1XOnXXfa+Y3b
9uSNkIsQByyge3RE3pOZUiWtHlF1GLXLRMN+rUjPE/PrA5QtI3tXp7kwOcVyidoR
1tjXsDBP75Rb+KLiSXeFtgWfHJ5m97VHcaQCprXazX12BUf6XVpk2aIExLjezrLq
P2bxpJGRoO+f9g+/m3nKCybx/mUM0um6rD/maMWcVBkLmsKYVkCQrOp+82Torayi
0459bnd4NfNiWSDAWa3Y+JD7iRKF1qQxy+A8nPLCO/KH+Pd5tRNcY7ZBYZzWj5VD
IWHm6SJ3nuTyl5QtE95rlrDXT92NXlRkhpNYi5tfXCa0QzPGri/cvvB8dzfZRTNv
Hnxg49JWzZOinSA7C3gRBRm5Sn3zGFGui+/Z54G9VvDldRim3+dyk3g3zQA+WPj+
MrcTHWhomkJ1Htbb8uU6BPlPON1UVd/29kRNohA7UI7UspPLLWDj0gHqXbREgC4o
RbZNS6Q8+a8TBDOVyjSj7r6j+aVEIowQOeCesaLhiuZNpItxErvUpFVtpzCr48qA
923QoIcBezuxTpUcinL/+16JRT7nh8LnOhkZVWQH01smlv/GrhAb0yHC5FzMhPsV
EqhSmSiX9BYTQzbmErKoeda/kZlUvoIHu/eMRIaB5WXcr5xZdMD3c0v/kjWwsjpo
X2a83IUaDdSO8Xc9jMJhz1qzp199GEHcwD60uDEmhzQUPXAYfteR7y+K/6+81lEX
0g9XevsDN5vVmnjMlRh/Cls8VxBp3GcRGb4OgQ+KMute9vHESXPT4sJsrE80dQ+5
OwCzIk+AntfZ7miIzKFD9UYqnHjDwGOgx0Qmil2L/xWmqLN62gpE3I4KK2MlEjbU
q0eYFG9Eh6g3H+S8KbmlveCYA94cd2FWEagSv1BiB6KVx/R9qFe5Ff4IspvV4gVk
vVvz8DS3PJENQzw3orcWR74C5qALX8VB3UNJSgrp2jMuiDSCiM2OKj7hpPa/v1NB
zRYyYhWTjFrl7FdKgQquDeKSIFpF7H1FHDjKydBNGHadHg5nZ8LFwYPri34g0JNU
UAE+OV38FcxIpx2CyCtNCYwL7wQw4P1MM5Sg7/6jCIuDcCSGlh7q6sTlKkvk7+xU
AU/lpnBE/FdYqvVTTU/OXt/N3WO9KY4Z8CjvQMGxm27B/6kxfwbTe+werOCEosIQ
IyxTBIb0B4KFfB9vgvwhbbqmAuDkLBHoi+m+k/Wu8cuICOhKBWYFITrPjv8d5QJd
sSGS+grGQStt0QtrxHsZLHtF4lV3wbpuCWgIH3oHZGCY6MneXFOYOchHjILQlT2W
fgcmb9va/+ad2nBaPp1y5q3fVeLnrDeZBKmOix1CgH5ZQSbHU8p1T7BO0KN0a7lJ
3VgEIdFghEuRPzZdNr7e4huykW7qcE5ZDffE1ug4kk9hoF56050s085YS/FBj9qu
tqqdrMqW8355uzICicJ/cSFayeJBmeGySZZuXwnegdKyYj/WeUw4RAcrUJPtJ+sv
FvnVIt4IHcTpCLemHJcRSvX/abz2SPSpsrk/dqMDbdMANbaLSXiSDfN1nbl0AAqx
47bbJ0zVbWrn3lGjQUxRJjzil60d3mHPFv83izgJnNrKvDuqB6kug1jAYpAgQQYo
dPjYGakWHtlJpxhbfhB0E7yxT0aTE//I3bY7EkdVGtMT80/4Zz1sbGkdzX+OK+XL
yJhT03p9ZdVXj3rLdNHdwp0ZmzMKfGcTY8RQ5rG25jUK4mD1MAcEMNO8/SSdeZax
cPwcNcdC8fELSC+RXzpt4ey2gt7E2wod/7ivBIhGFZoIv+YeEju0vkEHsslYPAhG
rHfeP5zfqi4sI5ycxhwoDoAstDwJNGr5k7+yGkZf3yA7abVcSqsr42vknYKIBQHw
h1TqfYnNoZHXroF2KDBbbbZE+Rp5vUWmE0FHoBYJjnz6f2OXJpjJh9RLq/SScpFm
1nSVQJHqbPH6U2ToA8ZBOpyd85Y9GdJwnlDxHjYBMDRygjCT7ph0Z/Xb7OTDDPaD
VTI3GHk4EJ2LvRmpeKD5dbFu+d8wAvM8+ypNpLDliScPDqfsKmjVLftnN44gRluD
twOO/vDXXeS0tj2KhbCCu/qd6nJ4zcsuQKLpgkvYsErPC2W39lzyFsi20wTSaPUN
DIaTDWTqpK5/WfTOO5OcKpNGw4awa9SUr3mQ/b08PXU2sH49cclCtAWa5IQl49Oi
UHqqHK1kiUDVBz7rtVxjE3FwfjtqlHJgBzxkZxoFaubkSYYdC89FA6P+NNAHVOW6
AnE1YL06NH3KWqFkcYeib4pgLYBg7ltva+/eN2U50i6wNrkOvNDQ44cQjJbwSPjr
QnbtGHwSaKOXeH4pDmChUDysYw5C54TqpVsbHKrHj/+N7cGMY3p3/5XrEGnDMYv5
NFQVSZiGyJxskewOfz8iHArfoMS2ZI/FLSFhYlE3sBJm73j9eltK20zxzGKdlidF
LaT7bbm03pPP7deqjYvm3Q3qe18sg4EI19U0nkyLQcxSn4lp27FYKtaRMDnry1V6
KddGSmILMCtOYuevD5Uv2+pRpuyWxLwLin/G5nmExEA2J7t/5lJiIMVRnY44NyKR
mR1z+s6bP1AAj8tSKged4PyOYbbTQOOhz6WLgAGMO5P/gbQufzYoX7Ste6kiQ9uU
KTO0/nRo3Gsr7/PQLJYHNvrt2OBZqpmcT1SXdPsvZH7ZDWuPSvwGEnng8e3ipAI8
5gJriJHIO42Ipof7YNmiGnTw2Ke2y3iyrcaDWUd0xYHKPjduh275fXqVIoL+ZJhr
s2lrwmexreEwe4pNNg8GOFli893p+NrYJJT7hnJcHYOz4HLVICCX8cN7ehvZ+iSl
usqUJ9O8cMYsiE5lj7bu2y+1rb8bUjJyi0psK4HNe0eC+HCAGnKQj1Nig+W6qy/b
v5WU422dvJHfl9/DMRmO2QTf4De2lCnYWaTUVJkjHNndxuQdJoGRo1tobDHZelx5
PzyeRlr8XfVkfxg+BCV5VPeW4dWfJhAD8sboGyOD6Qifde1N2WoZQxFsIp6GT5tZ
1f+FuODuQ+lQd9urKJom7/3SBGFZlte/0B+fah+GUuM5grKuZzz3jfQVDbZDALGj
TgH3sWW9JiOFhR3K0+oKZzycSVGomUn6GQ/Pfok9qxN/Cv/W7OSGCSVQMmc1BOX3
RJLuvbVb3qvPe9VmK+7cA1GPMfqcr3iE/tCZth+0vRWUT5vxLKPgHKYpspqG/Hqu
0aZMhglj6PiT+K2Is/k4KFdJkiO5ZNsMGpLIuv+Ono9A8KVTSnIUcRd6xzzujAxI
FTPXU2Y/TPCqZxA85/Ckh8AuS9Tco8KHebv4Gj7HcIi9Z2J+VV2lE+/apDFdcZu0
Mp3u6KVwJdcLGR9kVLDgk7Ht9JIT4dWNfIBeizIk2iRCJ0quJkm1z6E6frEc4KVn
mykuPMefsrP3/ME4MDLRuxHWNKq+UPmfuK1T5BZxtQu8u6vREed+gaNBdqcEv+s4
2Ns9ePbC9dMbtj6lZOkG+/SaqPedxO6Y10MellLQDmojy6xebWMZzLkd79JUq349
cAuJzNwxLvTlKAGW+60Im6pkVhZZRI8JGiv+ELy4c9CziUsYJH0+3DBvyI5XR00k
D1wLGn4n5/ZsknbiDfFgNhHawm8pyKhOaqivB4bnrNoenvCRlU8JLvIUvb06gy7z
KpYt9Udr9f/DPz5x4MKLN820rgAsG4JdzGcrWw1LDRHlo7Wlmgq6cgC0FXcSBMet
ei5IiTPVtw9rIrLP/aCs6zS29jkiqkAr3xLMQcQJWymloqEhICyCwuyniOX8Dfz5
7nL/RnJahhatNw3UBP5VFXRXzt+OpyNIyd84o+cpXDAU+pEWwQPA4pYbEWFWdZY9
TT8LJjp2PnpcYMOf8J4582PES4BSBnSokz7VKjOh6pLMpEjx2wFgin4soe0Z879k
Kj++IhBTwvzaGYd2PjKz64POCYy7eyFmeQMhs5899W2tOMfphLp4JIrv9qaGPBzs
PM7S7tJX6U6OkT3PPhstiE/RgbFEKPs9PiE3p4trDRMjfQVS364sHf/qTjYsJdR8
Bh4SyIHJ3NGkUh6RrQbS3k9KvOfsiHH06s95xDovbSLEu/ENCrik5TemhV/UWgXx
jSPMyY5mvcvygpQYFfRYy/nld1cr0PCRMB/QhJh286n/vrQXh4RwHFMTAl0c/4Y7
VyZ+NYelauKyrkYYftI4P6FxSg/tC7L+axQYotllfUjohDjBahu87KvbN/6ZIEGX
q4EK9P3kpULxj+SiqHU9EhXNrujEQhHqlcOJ3L+LZ2NLNwuuj/9VCgNKslGkCQrE
XwlNiHm0NORROgcUF4f43Hx/+sd1WMj4k6iTvgqwCiieeEXuvKX4nSwBh4hSJ67C
Rkcbp/SWeHbXT32jepPnDOGXKyc/Rd/vPD5VEjzXQnRR6CxSJSEm2eyivhns2xPl
kPGIRo5iksL9N7ZNYbQVu0q/664y0IeE4SfOabQoYHXBqZbgMMgr03Axali9p2a3
eUhQVlmrgCIS5nNuOC3KhW7wJ+i13RJVmB7p0+9tHRlgN8Lv28QlgqMgd8GpCMMd
WmJkcOJpQdGoNfr6jJzSSGVXV48FkAYcywh0SQKbIbF543N9ZVsVQVSgBQRlXJM+
HO00UqUGGtBg+FbSXkrdQ1LWbUwSDHTKXSXRXUF9V7zi8ttz4wwlrPhYtmExbWso
2Y10e83lnEPmNaiZWhrKmWlqaDJWhIJRn9C99xr7UkyyqKwUhIEEerov4tMWyhyT
UZjTVzg99sitt+T4OAaQ0tIcjKzEV+RvPRl8B1v1DwqPOrYfpugoBfr+IdOfQHk2
09EL6iq0D1syJYbv0CcRykNzKCedMgEM5s/5n+drXRvrXiPYvoD30qUKbt4PfbGS
ehcDNsuSMpz/nUAQs/EFKEe6Sur7SHa/qBj1j5RD/XhkAl9XwhFr2UFlgR90Zb9h
Vbo1iTbJPXGUKyKcRIRnx3C63JubuyRhfMTGdgxGYDkOjO6XUDZyctZjX2VCCZIA
NIqb7ArVUroMwc3o7P1BOwnWT5N5s6BQsZj0C8GW0kYVR9vHw/BRNl8ecQ3CheGC
Z8EDpc3xfnI0EGxJ8PXXGY0QtWte8gZbzTm8HCw3duMM1pm9cLKNOOUfWKr4G4i0
hliRPLkJSfihMefAB27mQN9pihUc8t94IuRr9ConehHhtYpuvF89YYdg5ftkdNfF
dHo+368kzZm14gV08//mbaGFQG4pGAFmzi/Nt0+5hefdiaJpyLVjotQksUhTc+IM
4b/2o5k92r+AYxi1IOfE6uOiAnjI8e1YczcqU74KreVvoebMyzj/0qQ+Fc8LeyP9
KkemXgjb2FUSkKWLojWzvrRqfeLDEJO0LR5tbxCYw5JT+lFkHXgFzgAQxViThrg2
+gxBuWPtuGSdRsSTp0cFwgH24glJH9hj+2U+gRgr3gmv7AvZtoXFquyaHizuQzlA
LfBhegJ41jju6JIQqQkVV7fyaLonSJwogemHU+NH6E8QekA32HTpsahFerJu3cHS
WtKeIkyrxrtPt3dyVIMY3WZO6XaAyu/OGH5Qnx1mmfLB9Pcpm9Vp1CYZYwcpc80B
84g3Ud630FOwgglXka7+71NjYw1jzEK+lyG388pQjd0jmfi3GS1EBmoJgCtauhZN
TZEsDPKMPUQBRzC3moO2jxkB7vCDls9LURkHBMGxRwlmtFUA5T36soWP7MrkEIf2
X6Iox4ZA7kEiiJ6HpxqFwyqjrCFrhpwvqp/58e8rgkd4VOR1LM3b4MxyPYbu6h54
QviXBys/a47+xr0kGPsxmb87ZsT40mtju/fILXXArxyGbfhfJdIMT4SSPa925m2T
pvXSVeqQuFDXRepJ6XZ3GTCDnfQjwusHFxpUJ86ayhMB3tx2BEhoaGBj9VdWyA6L
kT2Zg9/61q+50a9h0sqdBGuriN+CJekM5ZRDwyojdGpl3+r8KRQKUbYsCqJDYij6
6V7Getytz8ZF/2pxsZU4+d3lt8H6SNZ+LJBoi0LfDU9KH//h7qG9kE5hrqBKrWGG
iqhG31AdO3WyrrqZtBwLm9gdmifpxsqB+vYTvBuNcmtV39qGRGGdOdsw5Epvjhiw
MoLyzPvO/0c6+fw9sUGkxVNk167qgEKwx1jjkpmIYlFDiD2g6jFUpQExafWHvgB8
4/b03YCWaZ3VoAdGriWDRgvT4npnj3vGsvy7eRLq+vIGl64cQUD4RGsBEBSr8fke
jldlNmnCw+MXHmgZXEDaGPplqcT5IPfdAnoV+1QlmydBB5uTDG8Apl3IjaNsWv2B
6pZr9YkHi97UDdqMES86GkmEWWQR46S8u6xdzrz4glgTQVq1dXHrW91zho+Yegcc
fsHBuqM5VLAfzDMNnzQes4cODQL5oNUBXdaCHD8pgnQ8ZBDYYQmxBLFo2OiKxT8B
jlmixU0onQtQgp5QsfaEYjd/LUaE9GgwcpGb2OqjW8mUWWxrgo7kVfw3rtymGgZd
hmZPKNxfyQBkdCkPIbbv/JH1bPG9D6U1iGfADB5vFlx4TA7GfRFwwr8XQf9kLnPm
Hjc4ogCr9DuuXrLCJsrhL7DrOTePxX0r9Ca3m6c+39V/DMFn8z2uYwuy7le33FWZ
I7vwNzZXnARsabsTz9Nj5S2SCf9scdOMWALaLmrNmnCrmZhRbqe5imKaMjeFhRrc
rSQEbgSi5CR7x7cbaly6AuYS8ZDim1YHHkGR7YN/XVaUZKaxzdBRNP1dhKado67Z
FC1Ei3NgZA8kfy9Qt6bl+9Zf/Cg+gnqpNFAj+FaJ7nv8jHKhI11Fnvp2tbO8HLQQ
OfaJmn12rUZesIIDezSZ6fEmVpG7F+q/VVmp93npsn8xLJGPN9ep0jdvvY3tSDJz
WqrtE821hwd2b5a71ODDRfVyX+w5ZvVVcPagguda/7e6mZ2YnGathdktqJvl7DLL
BL334h3AdwwUfaPBvEirJmOl8QR4VhLInQVALUgKFXJv+kejiJ7y5OudUbM6NLIS
XcajL5uJxaVLHMT6k/xvClQT742IDoh5F7atsjoJp3mG59pA3HOHxcmhXmaAcOOW
B6mT6H4pgx0FC0IemEiF+9B39fNy1NndTwSa1cf6OuQ6Pby9/6C7QeR5JyPxVThk
w8/+qJkVq3xqFuRndNXLBEjG6swJm6qB386iQJ65Hpl05EAZ+ZYsFmlQr0nE3bca
cYCRlLHfd5UuLmhet5q6fQSNO5tYtt36+SBLZHgAcuYunJqLSM1G7GMPZxBk86S8
6mDdzPZy4bG4v6QwGFFnFLMJO0Oye3s/FMq2cnN2ys13JYny0yyy2BqLCF7g3WLn
O0XMXpA1tPfWIF4LDczCWUfmAyt2hK9BxHAj03MdmaAt3qG1gNnbQ4orF8Acf3bI
D7sFKbcTfHsLaG84iu27IfpGkOZrmmdjLUgAMSU6iOhXdq18Hs9/RiVtAip0Snnv
mRME0VjjbxxTc0YFGheC6TMgyQYMEzJDjvVr0hc36+L2p8VfLOHCT67VaRrxCzCX
ZyTdORy+F126ZzYLKWmLijBB9t3Gs2CBeUdv2quuciDKU858OzP+WZvEdfGa32nh
rAzJPa7eB+Y2zfE07+DUl/pgPX9Vs5ZRFTSQIgVX2wrBZ0RRoPKFNz/MFePMtl2J
fsVnfoLPhZZuBY5qxtGL9VgiyBPLuE8QZQ+gQzO2UyzkBhOk8ao7o08eiH20h9ku
B2+Vp/yMnwtw6dTq0Puu2tSkOMnXy5RuwM1RGTUkXBY7qi3jgei/wf51UI5YARDL
0hOC6gScGP2XoYGRXEsmTyR0jpeOjH/mai+u06U9VQujwJodKWzjgm3y8pP+HwYe
f2gBjhECWgAFiAI2PpVWJOrCJWfJ/yMfyaswuLUikSN0+5yTO2aKek5R6OGMUtzb
D5sG8WVFUzB96KHp84d/6peh56+idFIpjgyxXf8b6G/dsk03cdBRw0QYigi8PPHt
Y51iWDeUqcoQniwBU/7KxXgJVlSvjLFcm8iDDfzwJ68xN8DsJxdC5Lqd02JctCnv
H6nky8Jk6RLkqyCy4yQVxEMAwr1nj0UFx/0nytdEo0AmSeqLnCpG24R5y512Zfmr
yHu7JK9RwXDgxsWSgxSo5QKcNxlN317schLx6urZ+rqyWETQmowwwmWGKms1j+7Q
kU5F3e+KotB4ATizv9yFVO0OZrrqcJ8z+EBCzaAfI5o30vB/yLACM9LbUwI4lT7H
kF9OZqjIL6fiFEnWvtYOiRt1WhvCPAiULuzE0Xk/FkoDwyLnsIQdK2HVcu8kGbx8
I2givDP9jjiPEmirAT3osvDZ60Y9LJAXkiCVUKGGvL8vbpj9748XnC10es2yQ4sy
H87yWwQudCAoeN9XvhV1xQtN79NcxSG5PIDASajGM32dAXTAmFwmstiT213Bvztl
bAIVz+tCzCJVyu1PZtyNlZjmx8FX5H2idPSDgsFrCrwZkAeUehKBCPKAIpphY79R
kgIe0OneJAco6soh+03YRvYe6tlpLOjGLMSspH2QOgxE2Aq+Fz4YX7xlDZ1ryVU3
PK6eyBHcPMHtKue1ImHPmWz1v4/Bb2CE8drMf7wkdVp53dxSFil2b1TW4Hqdyd8W
5p0dfk/Y5nY+jvENR2biSPHU0mKW7+6R3EWJduJUkAJui6RAHC9phvh8byMnSAeh
8Mgg1L61rXuHXJ4evgnQm7jEav+hYZhpAvWfYZsl5AGVZMmHdPCtoAUKmp2mQUKi
wnXdJqVHyBRgsEhF1VfclMYkR10VPiDtAbOMf+0KqXYePD+1fIhUzle4KeQV7wk2
mQmzrq3GDx2DS99Rc5ugH6BAhVSuFbXMFj7uoNOTMTDALbsVoRrLSfgzwcwZOemm
0MR7kJHoa4VTarK9WRw46PtOPMnnWFtkkofmyWpRS4sRBMQoja7sck+Yzmrxdxey
3Wor68iQ/DrbF1lGfXZx0z4khmS5pqgrOb63Xy7B1l69iwPp2lIQflO8Dt8cKri3
j3ID/hdqQyuKLNI32AzhLVsMsKICJmGLovqQo1iO90qKn9kCvcGtLGSHwBT5O0Oa
PJBTxmCnpKRry6MdrX2OBYmiNKUFSLj/Idh+lYUnMvhuykslxaKr1LzuHoXBZp/S
w6VvanrB923GyzuF66UKjkNw3tZCVqM6NZ+LzkV7WIXHRLuq+C4ZJqEbsE5/9Ng+
eAt7EsiVBcc+fGx+4BbNV4pCXyfrnqRhO4/NSJuOsroP643bLopRUp1xvdMEMRrn
qtI7H0HMmBPd1lovnWMdRNUP0UEjQA89XJRfg4D2XcWqg196uJq0b6FxveijF0rl
NdNjttYEGIsNegogCc0tT/vSVrMGqGFuqmjOG6+1uZFNS8pyhg3uYkqSbpUpxtFg
F1ZRQKlxTmr3KiA4HoEWVAI80xf+curTcPzkRSlS09eVgRvRo9M97KLZqK6E0pUk
10wkaPIa0Ylp5l3AvaGvspnvyYgDUBXrLG8dgofnXSBCzcTM4CsFXNiuCCw76Dn4
9qE2hg6SBs69G2a2Xl0+eMli6m5iJmS2d1A1PBsBVsz0IkWc/zvDMbEEZuHktzFr
aoWhwuxGOT0lYgGI2IAPqJpQC0uvhq2ZlBFzXN7KCfBZa6x1hBGBe6WEvkmiuQ5q
jQWf3ftwBhI5vGxkH6aermnulzAqVx1WNDRObIHCtKqEhjAZK87Ekmvh7myA4x7H
fugOMEe9UEH7GzH81lioKLFmc38CvVvUogTyWlgkfz07XnUnmsO6Q6UCiPwohnzO
iqM6UAGH10aovTk/CS5GnIC1zscX3rhsEnpmBtlTIkr5rkHgzOrMI4yhyRahp4CU
XfhxCzmxrf2n9HxqPGb0nJL8gG6rI2dys3T60JiDhJ7usqsD73AUrFju98ifrTy4
18R74hLsyFxjWWk86TdKgifLPWJRokzFmziV2HOrBk97khhTrDHGrQbszGZHAfRa
46ujHbSlfVde54AcJ27rqx8aKmqNPKpfQ20YIzKxusB84qDec3KxpEUY19a/O/5D
8g/TlJtN99TmTyY7eRsJ2z3xtvH0w+L0XbqEMgznC0Qp+EqNy0pEXsCHD64rFiX4
O8m2lBMAWPB2NvF+IfrVSs0QqA8+QDfTB+cfW3ReQ8e1+yxLyptpZGhdqdm2dIP1
YaUbZKFVKUP7U4TlP5USaG9mkNcTKTBkuT6KWvD3CEupACHioB5g1wfxSnzvWMwy
8YMr6WOro4r60sqw51S5VdfUN4uZGTeQsT1PO8zM5u4yOHFdJHtLWKMdGOYjRMOA
xthlL5jWIgK7Owo4xXaa7MUYhDto7JN9rtwuYBEwo3hjNT6rcYWrq1n2NChJqYqk
bbtUrzdRxjyVh3B3GwkMLjyCtxSef9qlMtH0moz7rmFG9DN1UcX/XGZJgi9Mh5ut
PXWtJo8MwsIWI82LzmfGx5+Rc8kdA2yeBboJqqvJ8jAyL+fv2nDe7D5tn6U5a9JZ
tnhpSxVMa8srubvSMxxl1RLopBWY+ZaorYT8BCizkfaH/raLpAhGYfXRIzNZuxVh
f/4Sr2wP1xvRWrmmsbY26UJRqnZFxDINd8IKLfZg4FMbCTb2fekSj08k+skkvWso
y9Sd023vF147ThsqgXbvhdamyLXF+wqB4FpL6IiE0yLTI+HTj6rbrpVKKVUOjMlX
ZPmzIKfpfKVXXa2YKiEpuyM5GQS50So0W6chZQfrwSoVq/eJ7EiRMTdbz9MMe/nW
wQGbHQcAYgNS9gzLFgvAnXmt3AgefkhNeAZsFqnrGoPPZZX8CPY0NStQzH5VBD7u
vaR8HhtDkR0kQ8NqAXuwVQ6cdWjaCUlh3vUdEHIz7qInAGXGCzuWu7QZCiHxXsBD
b2t6PDyzL50/VWZDt+IrzNJBZ50jRpB1jPyWNnh98PSaqA4ScZS3hBNdgeB0jR0H
YNG8qjtP7TORqUE9sDWMct4Ys9BDsivEbJxQb7bxy9e+YFpLOPhnLlHoF/orJA1i
LBQSWrjRPZXdr5iWtxKyJdank3h4Z4QTvliqJD747uC0055EZOW1kC6CFwnXEaIT
hkObKO6D1P3+K3zd/sCJhxqwMAGjnzB/g+7+9Pl6qYDCvu6eSVvcV5/j8bUoIgNl
o25maA0n/0XpjDCea07wb32xgcOXevIOO0hdvRFrddauGD7cgSgyfy9TD9J7aDA1
yBT25D0ZuLYRqWH6Qf8CIauvetHWCpk8oj+DN2sdHGq9srxzB01VY2vXwhnXMzfK
fj1BrUUKZMCWJQsTCwSqgUhHxmkoh+vC4CR7HruA8mny7QVExju8LoUCNNdnAPx5
uAnyMtHgoGG2wN6uqmnXi1GPwmxs5419KUY24F0cmqYxISOIv5LVvxM5xwlRA4yc
91Y37yCZnkk4QeKCXcAqiTJZW0A647USo2gpatmCOTNAe/jlGvQTEB84koUqXK31
KJZgwNY9x6cRS7tbposjkwzQlqA2SaOntOVglVogXp/51sfr7pE/7kC0rtzF3QFP
Q8EmPrQHclv3jA2F702ANSHEjlHoG6wWBrxg2d2uXwV0baZ73IsQ+9XTDdoCULtZ
nYL5Jf7Mj+CajgQ3ObYedmnYY2Om42jydEPRGtR2ZDN9mSCKD6+eiyysLD0L+s+j
zgYaHkoDRMTvoAWYExhgv+3sU6LAsOu6j5BSIJdJ/fnICNHfYsOVXy2mjDXFIyPt
YrjGPQoY9RjIw7Zip5Jg3fBV+3PTNTELI4mFCoJzjRwXAzKop1hY0aKxJwjuKG9y
zQRrV3CZsRzMO7FE+0VMhPBpkUTsMt2KjrfnWB3fVlyBmXgLfV+YbQL5UVONXf1b
vnaHIgJ1YnEAIyaVKRLVp3faoNHdIyt/wiDXYfZxTAoUxVkpIesKrHdcSfLHeHey
nz1v1ZehoEryjwItyoC9mI7zMpwm/I1XEQeAiGCE9e2EF4H1Xwu37/b1gjj+qrKR
DabIRPliZSGt3/Fpxji4PA==
`pragma protect end_protected
