
module ALTCLKCTRL_IP (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
