// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:18 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vvxh0Z558MW4cvaFnRxBMMMPi+pFquIhL4GvjDtRmANKr/S8mupiOxBj81beD0jM
BbsoS4l+/9z60tnZpYSiB1l1Q8nmxDNCB1NFipWEeVOM+8RoY2v2wl3rvUqt14g+
PU75nnkbgaj7m/EKiPmy/O9o8vZCrK3KwNdzjjPcu98=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
Q+uzV0SO8Go6CzMaH4bMpo0Wn1ebOwO6oi6MPUCCXZOKJ9ME8Ax5vvnzjTcz5iyC
+tvweBasaWNruExrNHDoJSmlq8UjxyBvggbHDCJqEtEeax0Kg0SJd7j53hNi++EU
zmibwREW65d4idF5ruqFLLhJfGvC0fnaOXUWLCnE6Fv5HGW1gt4U5uV+agDrO3X2
TkHMO+IcthG484fyk4FEMrAOms6ikzsobGIz/CnbaIm79k6X6NjyTZPfj9icHDS4
/XGPGLnrEkTZtrGjYLDonaNNe8NpkFd6YELJiLdKqGVyJUH6EcYrr00ZsmslYrZy
1NVjF6DVzeCVC4fITjhO4iyTTxxRXANO/1/AR6dPo6L6LyXJSEIv2w5y0zqPCzOs
JCwssEW1ZWdb1pdT7G4eYhHwddK8pGoFQYSo6Rh6coieTzPv/UIcL4dy358kvWyS
gj3FU6kv4cFaZkvhFhP8xl2OgOY1HCN5xbIlkzb4scBBuMPYp9gjSkRo+lkrlh9R
iO0aV/Q0OZCesHttTmx6tJX/Hb0mwsEwf7ViQKM0CWg9KwLFrwl2xWJ3/evwYrep
FWG6wFV1cy7QY4m5Nkzq0WFh63ULwKs9P7oaUsAJcqOCIDU7nrU/0JFhU8y7+Vc2
EgDJ7mQQ5wSVhQX3dz4Fu4cout3tXjrP/WSXuY6Q7x4I9Gsa/ElwByv1h+zU7bqw
WFDyrrdkTgVm88im6BsWmiL82YwWdAi+NszVjb7SjJuL3tN1s0cWG4DlHhlMxAws
JyWBb/fE4njKlXr3+W8yX84+P6oGZEqIH1YEx8jWS0pE8qhOYoP/XNRC87VfGH3U
4gikrDOIzoDEWbFA/9LFKh0lTgkUW8HyZmApfcO0vuD9fs7D6xyJrxAH6FP0dbDq
sdoNieZU2WHQUuqJ+FHHcZ18aPcmNnD17kS83ma0UK8fMYHEbAVYqW2rgS7R76SO
AamiTZknj+iBSqk5iy539RyubvV67PpCEtsIdir0taG2z5bDKTJ/kkTPbw14hY28
1cVaotg/gritNYvbuutnpSWY5uu4XWAulXyXezXINTxzrR5/pKpvgYiiY0ul+4NW
r6AMUFs3YxjTI/SY8F9XBV5gL/QnwpC5giBouuAsWXBT+MRpk4+nJwvz2vtDKk66
h1gtcMFcELUaCEoe8ow8fF1/vTKNOaONddE4lfqnZV4GAYVhWaZtq+Kne3he8KmK
F19D4GFpb0Er5UhwHoS82TU74/4Mi+F+7jth/LlQR2s83ZOyVUlA9xL5EddHqO/p
zTkGEtRg2XXqR8DprwOxxZUx5S9Zk8pMhhS9t6RXxkm8a13adSfwjUgAJgM9hHuY
bwnw2KSGxDzkvb8nnSwFI0Fg76dL6ZgZclGKvX8CtYBfBKu4V9ZSVw+EuMYKqIGW
cBcE6fSeoHTDX/iN0+v8oij4ygdF/uM5UG9eJsCtpji69lDJbLLSDi/JWKrPQS6I
T/IEMbrSBuoIAg0j1uyITAWF/hHUvTb3JapFpuwQx0ju6/UGN8QAT3q6hvgnp3xW
gaXl14XVpjRrXH2DqmYOB+2qyJ0V5V25led0j/UUESWUjSVR1XJW0eW7UaAfvuwY
WUDaZQBoN2Ce5U1KqER5N2i+YphnQlzztDt03OhnskJ2k3GbLcGZgb5FALPhISFO
ysYlS77UDzlo0xMlvu/BaYzJMIp+08r5gwRQfNPeCqt34m3kd2/F4/vV/BLKSOg5
dIxWvpucpUPlA+pyR7SUJ1+M8bK4Ny7rpjcEhhBfz4ENcu7heXzR2n7P/2nOO0KW
NxdIgaDP+fbVn0aGyqE1svKkhxGcDreQWlsRJICKllKsmL72CifoMwpU6pW71V8f
s5D8tzhYBncfhvXaQIT+tMjafDb1TOVk3N+YW51ItxsFevwUfXvEQiWDc012RT72
Y2/fXWcSzONO58WfBjIeJzpVB/a8fIJRKm4tBdYidXW7p9UCwkUBlWhF/Pso7YTY
IfPM4otSFhJQzoD5GpwyTvZRLa2ZvdosC/XG4QrdqmZ8Kvt2jVx1UlL+FYLtDKDe
nsM2ZWiX3xyFqEbryJlCMHONuUvAVdbmBJzsS6iBWmG0TonBMSKu4DB97Tap8i7A
sw5gVXu1z8UaVfaubshs8iM5qauGr1rvhDSM4O1wbK7cJUQq3gKlrDXbHDoXIZ2J
PGEeZ498YhDb6z5Dy3agTTI9JNyQfHAmI40IaaQMY52kYASUbw74JDo1nJ06Olxw
li2fpfLXdSDpIGJJrmQzzhUc+Gm0HE6v2D8W8L4st6kff2WZ3AjLZp3SgsJU76ak
BY3T+k45azG7l7XrCk2UX2XuLAcS80pJ3JRiav2jQ9/7feTxbZnJl4cIuKfiXjBa
8c5B2JFmxuL1Uf/xapC3JfxvCFlibP0A9bcKpZYTBBnzb5UPa4rbquq82pOM1Xwq
6Sfr8v6IvrCG2XLuyBi+1NkK10AblfnM7MRgBjFc+vkALKH8AYi6SXaKI6edmcp3
G7HZz6ss15eRbRoLzaGEnPfov7AAW4nSQxx9VpFJn9L3MBi8ajTVaVWdOKJszqyY
qSz6452PoJR2oxP1JTlRuEuZ6o36z07HiUyk+Y41dcI0OiHQI76ApTHfjc8XxBaO
4wlXRaZLndxnf1OMaiHdJyYJLXieAKFkEKavA4LqHH5j+PKG7s3DppkeCujJIWje
n9iIpeb+fPjnSYz3kt2PAXTbHzv90NqsKKVuLjffQUoicCZG6Y8DHo1eQyGjCQae
N0OCXnG+Wqg2eNZC2mWfkdAGG0NU+9K7MLKBhSRYUenjKFbbU8HUOc+aGlsZ3ZyK
FlQuBl1D6RPD50cX+FegwKcP8inb0ImfiJ+71SW8M0kfxPfFwyIHDj2xa8oOjO/q
dUH2w7JwUuOgv3iQdWeHRT9cW7HtrQgyG/GzZ2xG8lXxKCyqYI6RDK8Y1BhDbUU9
dkS6kb83OUuOLPEk/WnHRliHrr9gO4OkOYuEf1iVFCJONEl1VJrZYwhg0nTxy14J
mOtYyApairiiBeIbskYq0hGURHavl0GEBJAVpQIohmD52oml/+FiFacZC+ZQtDao
DTjKfqUZeZMClSHpgESsE0AoL6OaBNdZ5E/8g0mvVSmzrvG/brP3JVuX3g7trnUZ
dznBWmG6LpZHpMdDV8pBHcM6cSdIbx3b+swwrmJFQvq6kfHjZGIXm05BQBMdtG9a
fT4BmdXSvd9CaaZ688UWPPY9Rj7eSUpFJhXjlr09vfEhX7gDllaqyAMG4qS1btu2
SwpDYW9uMJvWC1Lsg6djppWORAyznJuRLc13Y4hHOkOCACMmpsyDAlcpPZcgewIN
pNb6psp5oDTGpg0FEkkaXeAAHj9efw1N0nBu516RY57+6uIHLTH4+3DsYc2vqokh
vHCY+5+D2Z8VQeG5jc3zRJygQjveiadjWNMH1IjkuGggLoF6pDpK9EdiSA9JTH38
39P+qNzdytyZW6uUokNxKGRnGzZN4NNkTQr7Dwa4th4mX+EeGjH0UsJvAUvR2T4v
5Lr0SV8tXSIbXIIltWaKSIqz284+c8flq4TJtHfiIhEBHCcHqwf+dlFeG+xr1e7t
JArtrSIr51kI6AOaSE3t00Cpx/F9SUqGduzreIaxNm+CDEVMnCANiDBWcex9brlY
1NdsK1SKByWooL24SLf8UKe7hm7LkCQalVOo8ZH2qzo2B16Y2B5lrB9yAzrLEkYj
jScGD7JAa0M4/boCeTEZr4XZpka4wkXMWD/KmE/z4/Jp9vIKvmeAQOViGDUoS7cI
a1RQUIbk8gvufs84+q51QmuY2BsnlcWPiNnW5mDx4+L2d4F7byXOnAhFyvkt13ky
Fc53Y7sTEeSkYGncWwUSSBw+NaX8QJfXXoR1oySAlEI/YskgAL7z8fN4JV2t+mom
uwy1U4kUp+lN6MUvi7gbjT2pqk6sLvZnUzYfQ2I92Fq6jSI6fECms2UYBmSOgMsO
upl2v36DSD19XNU4mf3mYIIq4/688y6+NdR8yxFKfJXhyIOfbJ5JTacOm6qsESbe
y+J0LJL6HgkPxK0596Z4rptDGqZ+uZVtFk9pW5EwIbBi90BXiea8Xc/7FVj6HO7L
ZnFnTHaxENQOT6hVG4M6FZ/r1XkEeC4EjUb0lWlIALQRYSBfXCOVKzbA+iZomUk2
Tb3kghwS8ZSZ5PkpOMYH4JARnzxt6MSdmryIbNATLT5L1HNxNAmnLqRgoWF33eaO
jKJUiFy+UpNWUI6unn6FI/jDghd1+8vfp6WRvdOdsJiapnXTgQieI3ZrECC8MgkT
fOJIXXWZd5t1t1NwQTH5zfGlcV5M8L7hr2Y0Sb2SGiQsDzVrSE0ncF1ptSIOGMb3
OGvzAr3x3o3DcmJxEpVkjSSqvHf95Arkcr4q2TqTpVbGHCOi1YHp1o+mzQI4fKui
OJBqW9Xf4YVXomKYAPhM39N1DZKScxcjGnIqz0WMJrVwkso1xVxRApy1RQjul6A9
kHCzdj3iiYgaitmnnRtZb8ER6gpne/pUDf4RbSjMLuH1VV4ia4kGdctlu2gMVtKW
krcAJ+TugQmbjWTCMggavDhXwz4pLpSV2oEcUI539QOlMn3AjVyOSiY+fd9ta2gI
X5JVL1PhVPkU0G6wN71xLx0Kel8gieuTPCuDfFCmH8EJkQthw/YUL7UefdAWMyNa
b3APdgsuwo36OKDfuuwF+z618KxWL1d6hiW7tuN960oibExtMEng4hKie/GCHbgf
YVDJAKHxtrhkhqZegiz0FxngNzEqRf1LpxvLeC9AWcH9bWCqEtqLdiJxDdK2tyyP
mkSKkZfylgCl9Ih0Er13Jn+Y6N+U7hu2O0g3w32zs3aAsrpmzDxPF6I7cZ8tvDD6
jpbrbx0B0/OwFq8kEuirdfAyMEwXIk7/IUU8dk+ZKvzLDu7UHVv9FEUA+FOhq92C
3ypEBa2TZi9OBqzVfbx58FA1jN+Jjy7DczHG+oLE5sKHv26cXl4bhcCipRj/f209
Q5IVWCbcSMChaLJMV0if2kgnJj/XwBZirhJBuFUHBSO+G4gXSAIuWKQVjNC+bkKP
v0t8qNj/Ax0AIS5MPf8skdIHnXx8SXVAsnfoPvKjljcvCrSyqrszky7UcO/nZ0ZV
JYnhcvEZyFJ4aGMX9duhov2UYJs7e7lri+CY798HnbuhM6OSLOg9e74gA9X9UeO+
GksQvzDdtac2BCVfHOXScmOS4Jv3U1euoFRYH6VzQpXdKZvJOGBywuq+QhTIybbD
OeKcnslAm6JdqJ2V+okGYyFirqFbgH4Gn2UwhrSn+GWEZHHoHVgK+XfJ8D5koVor
9qM5XY7Fj4n7Vhf95gmlOrqVppRmFEkRPpNNYq+lpSNB2EmfI4d0M8UMuAPWQ88f
k2bGiaPaKljOcwSBSfzlUcGtMYl6PFCASIs+LFWze+EdN2fhU2LXwRzTPekjehYe
xFrmKKcVAqYnfiSXXqMNVIlqBt53TES6yudLn0TYUUq6pxLGp4fs4/rxjkWFcL2N
7nZXnfyPUVBJh0aG2yKsc9i04Xk1NuLCXNZYTHSv2SC9k2mKKc0eSFQfrE1dsKih
4/kjSbaxd587GWqEg8ZJI+fDIG1l0y/pAp5JvrRmtUHkV/+bUDlSf5HxqD8WUj2s
mEVv/oS6gZWbuoxTm13Erdcz5rPNz/Fx0JaHz4jU1BXyMx6fMXA0SXz4Ve/xXqE+
L67kiFt3FOeSLfo29lg+GuPZytmXehxcRYDXVTVBqPjK9WscotPbD2XIlsOfJFRL
WNierdCXQLfJL3/RSQ58tVIZQuDX0Hm+nq5QRb+vZ8kokzvnA6frwBiJWoH2UeTP
GiFypUF/xdEuuW2I92Uj/rNtq7ExBxoWzvbo70dITbYhbUrtMYa/bm6404fQrF//
2zbhObueZWnz2WJ8BUeurwclRUFBrn4bGydspby7WplgZtQtsdVGowhsiZ/FHmld
pvMSxneSn1+5ja1Iltim+7sd80PQydF0ievO81sT4LzmGDro3hMsP1EtzpGSY58I
tCqB+DT0bi+ufQoLEmZQJmfW7vjgBGwELdArrPPJPnC49D9PmORVK0fOsUA8Fbiz
7BsSTw+BSbfpSRt4F4soXCfEwm9sDAxtDDwnC6g9xEYrnAPSOJuFq7CCmLqauSTh
7ZZDuBNjW2x3tU4NPObQsVXLzscTX0Vnu/q+ArUZTuW9HTvf8wrL+m7Qtw21xYcI
qV5olTyy3dZbJZbWva5nFBdLR/cnIDm0VPNm+ScVYJlH9injXMseE9ZsCFXecyUo
9bUNxMX9bC9RWSs2o61W2Y/ZvNKNd/gLfZMXu4pt0az6vj2zst0+ojUCSCTt8qhr
wlU0qyr+tsL3ZR5Fyr9T6yNFSZanfNh9OCpbWzR0zMyXJ2jEnCpClo4WN6/kg3GP
z39vciN3MH+yy1fARL5qTaZ7GlgPzySx32N6SnpGMZssuk1XC3xQYPtlv67T6ZfA
dHbN6BaHy3LOtGApcAwJJB+6TAc/cE8MDbJ+2WEp1q+PxTPENXLXGh5yfCWmTd9y
Xh/G6TpVnwJ5SkoPetG31AIWxxiSuXH5ILx9vcnznIoz8B49GtKaYnvtJoT2KyQ8
ENLAx2GW+0jqm5UB2pH10fXAZJjxbVIJC0MUZ2fFkUIVBnGYSv+7WVR/YPHeACyP
jM4VdtVQu29H/pfTUF0JrgpgeBUQUrVuZ+2TngZYvGsKXInXCsucfH2qTUFhHD7N
NmvhmuunuFIGWQrGDzKPeONOxsYkhO5pVLGJ/i5K9cAPvzXjcQb6upnlaen3uif6
iwq6G5NUoxz/Kft3frPvxOeSCi3n5USNrDihVnG4xIUeRU9NeTRMDRGT/cBXpGVl
HLNQx/W89KJozDoY98gFRRoJJAysNkRDhKtdEGo2AJ7w8Us2seYz5t4qCJVbrARL
AwpSPLm3HLjQKyi+RbHrRynlcRtZbMbvRZ63OD0gR6YmIzJiPpDoZUHrLOG5JNbA
jE8kl1XVHs3bu9ZdfcUjHP8cZhSh7v4r5ZqFZyBQuks/7PhS006B68xd0oswqEf9
E9XHxq3gVGL+NdaWg1wX0IVYRfxT9UYuFSUPC430EtCLjLJ1QhABBlHBFFwELH4V
gPGvg7gQwR0N+BsQIArm3Dl7MtoAvDU6J/6vENLQ8wpumLIljLQ42A7Z9JrnrKaE
oFei+QVo0LU97U4c2PqJg7zUmsynMenFJbUW5QoVziQ3o58ZKGAZ6yabWIN472ZD
aX/XFQScCwkYRqVwpZmdwqRLbjF8U0KyUqFwGRPYUVTj5CUYh+ptE6aOh9z6wreG
sLie+Qje+edfq8CIMzT6UaRFq2Eu8+niI2tNvCqNf2InkMvXhu9eJPqnD3xJSLYM
Y9aaq1hrD91Mlu00eNeS/gElIpznvkREu/f/sXzufCuBiTqOKknSiczJCzlUoic6
ENu1IEsfZFOi4TErlDjlF+nMoAKYnEvOWuB49OjAw8wS4ruq+lzclT68Dc9PXGQr
LOwh3WrKuvheC7KNQ2HCQyHHvPR0TXzVuzvrKimjZm/Nhe4QHyOJeIbxVpWDwQz/
qxTjV2PsSrsQeJ+2zBfi5IG8qeHPP2gUVNDO7jUuntpxebshIG6m2aLCCrVkO9Z9
WYhZStL8l2blBlgCRGd5Kdig7bFos4+hKXFxLUZ1J/QxrMevQYeaHt0RMTBg+RFV
fy8JVR6ABLBDUTheYFsP8Ddda+58v91Q1nG2Pu4xwcA=
`pragma protect end_protected
