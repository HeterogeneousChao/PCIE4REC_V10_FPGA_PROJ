// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:17 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K3CgCawrbDHhagh3ElRh1Kogx40FH7yVpqcPqQgbwzuBj8iv+w6YjM5ruGLqK4vj
gYtk4CxSKk2lv3sOHK8RIJiCwtxM6dbOPPSB1okKWYbQqv9Ecty/azAa+g1cbu+8
VLDLNhkYBofisyj/vP78YKHeclAzXgI280GQN4KqUQY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8160)
L+FnuBYPMcLknFGGuP5YvkLDbGiNtbmKm7SP3k9jtyeaMT2+yOqMWsRJfa6iO+jg
zrqgVVEFe2f1+WlsxEVV3J/lP/1Fudbsu4cBzvY6TCXQPXQDgKT11ma1D+nwQgE+
JE/FwiuRlsbJwUGCybhCIXpb26dFmsM+3G2cgx0T1cZrs1O7lcQ0Vf9+ZZW4DSr9
MjX7MEUaXAw9s366RMjlpMUNzkezcY/YlQmYAPrOexGeQ22tVLW9A+pcxYgoDaJ0
YdJKo7RAap7Y2LHSpXkL1KsgoVFSWe+xHkIo5esEap0+UXvez/hQ7aFIY/pjICue
uW4fruHyMxkmGNEqwmLhVk95GHAuTKst7Po0guKYj7ZwoBWBGjTT/LyHLpZ5c8LN
dhI1v+lj/cVx2zK1LXNTh84idjFnTs0aOD0aYTxMi+D5GO6zYUgKHTo/anoP/41h
SN85i/5wVp7hQ8ywIY5ks15nGA67yd6U9hHW9xenfQZgTUQeUc9i+vtU1BTsuR5/
h3A8wxXe77cpdqbCCF3gotRluinYcOg25qpPVpDCLHEC2nwGJ3wMjTjK/Vlj2bdN
WcsrzrLAuXUV5X4w5QcR+AY466gMUoTI2muBIpyywEgNdclxW1WMP4s7gy6Q8xVU
LDd1bHIWQzhltoIB/490L7gy3+rYhgCX4EV2YkbiFF9heRbBZRrdYMAj48EaKtUs
JZWvIBhtSwgBpXonrFxf84F3o4IoZ3Ds52p/7XHCgLE3Ktj88Qk2NTqzYA5AyDSL
kpho/AtopAR4euhiAkjqb/YTntoyoUcHqhmG+b+VPadMIsuQ/M1zOdjmgfS9wZnp
CTWNdemH8zATse2//W4TKHRwKCiP547czJBJJDp4bQA4WgD0B9ANuL2Jr3Gg5MuX
/atiNlp0vPOIwKp27B0M1Oon2p/Bcx30QsLtiwmb2FxAHwRXcNWwMybZRfhiXuIw
tE1F3ZAZty4f2HgnsZ12Bx8qHBe1HQk093wm/FQbxskUq2D35KQPstQ9b5jFiID4
s2Msb7eVnQp/ewIRBz3ccBCEMn2m5L6uk94UBtJj7PxW8CAz45WE+SLW2ZU0J0am
99SGJLHBkz0uODSf2D++ywKNS4Fkl2sHV0+3yZ2jKZHg5vw7gMQq9u78ZBP7kZcQ
+zUI3evkdD6o9DCS5lf7yXAA+/3EeHyhJunrWXMO/NnQwvw8cUL5J+tcVe7P19KL
/yjkKV5RXdXAcDlmyOLw5MCwS3GiLeZE/L4sZnIMhngr2wQIABAB1ZGuAtMuQSjG
/V8iV1taXh7MaSigu7Ur5geXuQh3e8XsC386sOSo/XcJdE3SIpXC6uhT+TZyyxCa
1ziaKBOh1//4I+DiivYd8Ye2lawflpzQ1ujCHQlOh+4SWeCpxz8TqcMK6W00j1eF
1Je/RBl/NkvtsXW4yKSe0esmraCQmb5sR8iP7QqXQcPT4D822AaB7hfhDO/gMflO
WbDONlFXPlZmX7i/NYTPmp1qnyO3KC8wDQtm6L3W726qPuZMq8ZkY6970O7UG+WM
KRbvy/pcZTgrZ+KK1vOIstBd+aj36E3+bnGzx8QY6Y6z/Rj0e/ONjDKIKkHIphyZ
osKBd5FNv5CXyjIJQwTWzcYWeybKIKxWLOx6B9fOF3dz2BzFzeJpmvzy+fvXjjDe
lMuosBa7EwdTGOCjL042SByRqt+yXKsoux6CPy70nR1BzxJ9dzekcNHGNc3BSrws
QiF7sEih9SWcm60J5josWiU81DL6IA8kRZKrkn681jDzlZNfrP+g5mWF+NjgDZf7
bNZvZB6DtHSVXKhDbgcUBi+U65GqhQRAtUgLpgnv8dj8Fjc+L2Q2IpgY6yBNOsZL
41QPXj0aPzmtsG8mshW8kbNFpVVfAU7oJvmaTeoyb3zyegv9pyebYhGJGI4qjmjm
8PyHlIbWghJcDa+QhO1B1wU4pd6PH7mWNYttZTgIcx81WK02xIWTln+h8v1KyHYB
VGh/YmLKaU8pHhOZbcz8KoPtrQJCF+syy51P47NFdqNudRS80R8pvDJ4ffMWDzd9
i9cCW9CCugpJ++mEh5gRY1s9AEmucNNmkZ2Gq7D6SDs+lfjqfc8MIS/LOJaAZrIy
vagD99EFBcf74/nwKCuCYQ4RH1FVWVr93i5b9IPAgoOskJocQcMjiOYdHyDADrwf
LJyG66K034RC/DHNUuHUnO4q8Cm2BylW++gTxmhbhVdkYULB/dwMAk90AxjhlNJ6
8IDNR97ISPoILxxptjfLPvZKn16I2jyR/w892p8l1GWCDnkE5inIsQtUnFs6NJPf
PKMZC6OJ+RS5/w5KfnDtGqHnfAe04eUNdgHRKtllelU9vYYzCyfMY8gEib1Oz1zJ
79YVtu/6n4l4Cw6P5d7udoW4lbtyZahj5fidRqshLifpE9dFLpl7ltfewR3OvjPl
es/rshgIpNtUn4fFc+2520flubgyFSDLIRARkJlEPKBhVd99g+vN9I7lI4LgzpSF
jW5f/YgSxscfRNC/Ad+3jrCoJRaW4cS6Evc99VfShFLM79Pwi+IdYxt1PvOmqUfs
rknSHGMTUygNy9U2KJyo25l/et+IICRRNSb4I+uSD79ylhoP/UJHgieZxj1zKuam
UuGvmmIx/emins/Zdkh0WH4BQFGgdWZ8wcdbxYfv7CWU7KjPuRSGF0pS2wtTd/ri
1FBzregeIrV+KnIv3LGjg7x8ah09f1H4YSmVtH/DKvh1L1pSuw8++1k+PcPKRE9+
ucPWuBF9dmj4Mj7y6Em1kAsufwmINe+mUgbiggDi6PN+q3M8kpVXN4gaAl4nahpa
rP8lzfY2FcCSDlpQjVCh4gUCzdr5btDgR3thIVBnloeRRZiWuhGQeriFXinMscB6
j8DTSAb4K8rjdaGNBAjaOSMv/iBstnlRe0Ldj5y1V//k0+S6aieDU4RfE5ft9q00
1yBwINVEve7W7wzpdO8ZpEOMwX4wfuCHiMXKFxpJsZ08Z+oo8FiuOBf9BjiPkhxP
zy9k6ZCCTmR7B76ut/HAVH0r5XeEU0U3CVSUx7KYqolHjAzNX3uo3F9+3B7msJKX
JYYSmVQlbzwlMj45fR9A+xeLJKukIgikifqOwG4+R+sAGvsPMTBG1XfgeUKOGDkg
y6O8bcHFfYSR64ssnnAQNTZy99i7EZG2QS5OB+9gRoNExO3hed757qjd8E0uv9b8
SaRqmrvgxCxjuEuMncSgrB8orIo2VbyfmQj56Lh9rIQP5TyTQeWbb9bmc9vF3GMb
yBpwJ+fd3DHxRBf1XDitKh8kWysXEtn8V7mz3OmLzUMyWN8d4r6xriYfirv6RGJG
FQc4wn74ryUl5PtSNmybScf0Wg8Xr9++0N2Vn1sWR2OiOikzLzYLkx2AOyksYnoX
kJz5N5clCkx41LXEcs22LoZ8ONNFAr4iEZMpjQP45/mlqtVWgkISL7aQjgHsmj5n
nQOJeyJOhjU5HZWA7Uh1bIGGz42pCxDZwxndjhR8MD9/wBKcgTUm3NX6YBQAmmE5
/qCz7i3D8imD1eR+UeLViK8s3cJB2TsNXgVW8u4tabmLb5XhzC3ApGBgqUhfK9Mx
6F3mLJ9ByoJbq3Yivt9ASfRSIJUGonz2vkEGDjxSL6R/1uE28qEyf6jE07t2otQO
ULJuTZHqDwczirxJIC/Ky5w8SAwGy5/hlWPzWk7bXxRUc9ONDaJMtHqGhmw0khe9
EJDC+WMlkrSUuA4n2/6RwBHtdH1/yerMTj0IEEMO8IIZD5qjEVFFBmWh2Pt/3pjQ
ISJFMQyvwQtzvbmVN97lMzGENu8tZNtNnrOITLB1+s1ucTWF9pOcZyczegq/vJGp
Z2akcXhxnMLYTbdgByz0/OuY8grdE4Lp2xOAbJdvaAHYwugNfa0JYjVWSk4JHEhF
s3VE5zHVAtTciQu4+hxqF0JY6vDT6eCMLjBYgD7jHk4jV9D8i7f4Bfi0COhM3ABW
sjHfaNMseDLMSck0uAmdlbhZuRQa+7zb20Del602HJU91ahoP+GIkiSAoFCFDSfS
Uji9Act1VmfRvMX87pdF2Syce1odqEbJcJ8T2Zc3G8ypsHNydRuf5N/lFxVUGb2+
Ac96Vgj1tQUannIBT/yUxR3ZehmZUTTMCZb0yBEU2F9azYRupLPKN2IajvH2GYzJ
livoHGtcvwZODnROSLdjF5+5mLwPZmtcuV2OlH36tuuGkyvPtQcja+C6HLsjkqDR
JYJ6dHHJ1MlpRAPIx2HOOUI/fpqoqGn3+7WkGiULZU0xLz4qrm2QnsEeHSbTpfSY
y3RXvg0ennY7tBRcb0qBrmycjcojIH7xuSIoJtHE4aiKff0w2I65s/X7SBVdEFgr
G1epxLp9GyxQ6U2mtElB1iOOtGB42PLQQZTachowF+4ndZhEUl/T6tN04UMsGget
dBrX6Zzi1+7DIXxL7k54kkBv1G00DECoghKgVLVNPiyfMRf6D0j3pRO71VHZ9Uwt
8aVVEJcemg/kmd6Tn5dTXQJIWzq1KogReHv20oirzGCs6/GEa6pjJ3XWRF868z9C
AYZt+gh3+P9fSiRr6whw1cuVSLuvuE0lTpc5ZxoZ43nyxvoeQ+UH8ZoTMPnBzknr
ROQTyGKERHP54ue36Eb6Gsb4O5pAuQ6E+tkEyjXO+35CxhzngbBXb8F4pixGmo4u
MNz/2/nw9oLeJ1m3lRas6InHzXlmVM1q82t+CAdws+ibZxlTsxNuO8Hndwcm6I+a
CEncZlIOfdyY+AQPcE1n65YH+jOwtQO1vObxow5LlfpTTc1fOO3INaOV+mm36b1K
Vo5ockQJCBGcm8Bo+1mnLCpqn1mllxfIVJLxlIob/spxF3UxsoAElVfAa7wDWWia
OWVZw0r6fNqOf2YVGbNCF62smcLEsmLBhhNHNe0mF56mSODFGEf4cyLfD+l/urLL
sIuM6btjzmFqdJpOwfNPuEqxzMpYlcWwBn2aGpDutWXZ+fk54ZY/d9sJlzE1hqDb
47n/+1kX3Egie9SRq+Wb7VuUfIJfiplFBQPqXBPzROrBHcKmxRZIbKrSMt4sWcdH
e9VYl1m+46m9vxXeP+hTeWGLZLACpiZdN1tUMcib/tbu7bFaxIUZ5NWXG7JqbDMu
r5G67X+FmUplHey9/LbcBLKdA7vDQJD8mtjT6rtazbSa+C7jQCigrO8GtyOI8FwO
SA8CfZIjGYmCJw+JhQ0XmG7vPkun89elFl3f6R9wLXum2HHESkGwLH9wg6BvLH12
NguVsHBUAthiC8DBQekgBQYfxLNP5+j61o/KoqyoxH45BCbY7ulcqHuR3KKtmdT0
CP323LjKRaqx6BijG3N0YZSy5qclanwvWNtHvJ0/F1W5eTWzsIXh7Gu9//6KWmBR
dqVIIkpgCY8L/KRDAeGCcmhkI+ZYDkGmp2xL0bYW8M4bZlaeSiJISH9dP2MNk8dJ
u3/UtOZdCJ2hvSVroAsLAR96FaNRYv3uMcQ9cZLpmOHvai/OtwkvnIhhSwe7yKhx
XWbNA7AW2odL6wp/EcrQlAYzJrHI5l33Pgq0tXHynUcxqUe53iw7GfDx19Hzhean
b0pA9jHgT4cLZi/QHYuUFD4QiCslUjjAKZ6sK1ZC31QxlSHc0sXZTZurOLy7MKgl
grKmOj7meelQCAugS8vZbIgjmcsz5Pfe+F0H1xeXjhB4WXqEuf1BLffjVX3E3GOw
EBvx0ATWXVxEG00wVDvTqMTTsiyGltx4qAo6O0dgRiw3X3+AMFwiq2mTHSadeElH
+yaBLPVrRvLkOoK3GP/5Xz5Aje4U8PodEWTnFfWbFt8uSk3v1VgJOS9JbFWN1sld
2vv3hWek1HYLj5YcRKM/qbOq+HYU3V+fj8f6QG7Bs1d8TtrQcljC0Qq+W/ufCQZN
vaaRXfNzBbLard4DF8zs7UXuKXiG+sobfcQIaExgtCMm0sy9uIr51HVLZ0TA3YOT
YsV/Ci4LzWvJtaxA6lPPSgZSDg776OWFKas9vrKsHEDOjCb2qTSwnZ+ngm4yOtxL
QX3YvxbdqoIaSP+3IytUPZVVM/M+Mp481i1FOUIAkm+wsxM17LIDcXZ2JMBv0oAQ
FLiSCWM4rDq7NDO7+UG75rIzZRLxmaNz0GGfcgqSdvM+5WZnuBXxXYoIhqu75sAV
sMbeUP7vti0Zrqtn/+sn1rrFs6JPwcH5gg1V1ahoycL26PtQpiSt1pIBpVTDrQ6+
AvwZ+eJkJkf1eSAODWhlFklGtBvz0bheSyqQd8YJ7RunFGl5+RTqAufH7SwtCmK0
z2JhoLSbBc+uOr7BeosZi2rTxjriqdLONpHulPlnTWYmEg59f8Xv0+Uwba5RtOBU
AfU7cu/PNDfdz7Dn0N19Dfxxgp1EgADoH8Yw+yb++QtA5d0r1DVlyfzcvnjxhU2z
est67le52wnE8k0HFPf8ikM0Xt7Tohk+1AcDav+pMzko4PkTpGuVrdtrR+/wbiml
Fg7yT0RM/ofBxcj8bybCM3QVakZaZ49V41jEen1PeqVNEg/haBgaiZHnXGINSLKn
vXZd9AKZPikyh4ym3p0xT3SetI2ndgM5NwGOpQrv+zHphj+ZqUkRg+g6BvYevOKe
YrNWoCyQP8TjKLi+aFGSTUPlOnuESbroXgbnRfLlVYk48dKYYicIL8JBoksbdZnb
ICHMZdlwGAJM3DAgT9WL5QyCViVUvYrht0taYyWw4SgAieYPU99f/XJwEFMJB+By
F39asFtxL8nG19iBf++FH1cpBn6yZdLHyuUz7Upjh8FBRyMWi2fLmX8ksZud8NmI
cg6pPCU0Zrh0+fteY/REAmP70iTLPRBiGkKuOLJmHw6hIzKY9XWKZNXVIydbTVYp
0P1/9XZiAbymbgL2koh9v8O7hMkJoPUkVTNK16xv9KwGz//q/ZNvjItdHXV8B63l
KwizsntGopt2tdV5FB/hA1JzHIAmnaxiiRbkh69rGYKCaklh70c2WlGhT1kI4i7/
hJFRH2C8H8+Ja0N+oTUysDJ/9zD08hiUbK2QONVSOGwWI8gUsiAxRzPPAxmTgdbd
wdZpZaKBkCu7cj8luIu/72E42+ynRkfZz5Vs4ChyqBMfzhCxnQN16BlYxu1LbBlB
m2YpOB+oJi4thOQyxtRCTi6ETzCdKewv9fSK1D6dD//orTzyVTegLWVXYreavjjK
cb26z260mtG8uSu3ko4j1iucObeOM9Lt4xm07V3+4UeImcBdM6oBuRA16rjnpjcX
Ofk/Vtl3lLx8Jx7b5dWKDkhsxAx0Nimcq3qDwNlphxnUwsFf8DT57juB0T7DnkWe
A0CH9LKFszeJr8jx5Q5c0ESGFixtAasRS8U9aT1itzajoLlaWYvOCqfEDT1yudjm
AqvDcxOWriV9g5fRZYw72autnLRqqB+MqR6nFpgOBa19Onp93V99CXJ0IAQKrasO
9j3JR5pc6iLHWRZnlyhewClG+aBOzfsMAYkKsqjRjkUiAVRbj905dYZc6MluJosY
aUkdqm4VfOUlkF67cizVTRpJhqH8Z5Qn1SA64QgTs9umaHl3VUnHqMkeeOwCpzim
soiWoAA7I9IivNrdLD03AS7b4svU//bR8ERhG7P+RU/qePXKMrkCZvakc25QQFmN
3xD9IpY0jXcAQObm6l6EK8rEOxbL7tbFJRa7QstcCPxUt0wDgMKdL3mRtMLTMNDI
Cob92/DB4jHRaHQ76VaaA5dVd51UloFifQBHIPkuWjhLRinyWFzZFi0rvdjxwaSd
BzXj9AkJn6qrcR13CSxB5LWEPflF0zXAxgzhP2jKMpszsCJU50jDj4Uy2U2pVH0n
RoZS/8DqtdiQDPmD3brR5c5WnHmMhacbb/gXTwpEXkDcv3LSldHguSiaYTybMfju
QYMf10rp4/Enkb90InYhSDQSXAKaiCgOFRNTER2ytwNsP8FfrQI4GRJjyakVQDfz
Cq1Qt3A0dMltUKdso8O1QMfIILXLR0vfrLcMA8n/x7im6YyVYFrxD/QOr3PIYLW7
h5lHsKmyrTjSNrMLl/sUyKptSSDjcZpze0u4DMIey85KSoigs113r3jv/yj/148o
P/IzXiGZGsgHUMVCmRvC7NV1F9rUuF3xByLS/J5sDpPxD1bvmwi9OLtEtZiPCax9
BeF+zCb4y1TW7hHO0K2biOZ3cyE9X69OU31y1NNv0hiwOOUBjd9CIHkrlodStkAB
9A8Ru/0WgQlvhL7dlsabjyaCJrDb/ESvVv99MG5KeRqAIHFq5xyXEfMWxDVaIg72
93xRrMau9chS3x8LkpXz38aD/sLYV2vKiyh8WyLTt5bJ7EoTBdzts/RFYb0xp0ER
j9HXoSznSIjIU1LEvY0E3JcnmHzgOxoeIsysu7xmO0sTszNb4BjExMHjWQrPrF7B
LrA4mKkTP+Wcr/9RygGbbJ77E6d0uiWVeKcCJEDiCXfKyS3xi1gg0h0waxSvhzCH
Vz8WdcQJ35dEpQOoaC/nyyGWdHiTlj5GJbnWt+yGlbr/1uSa5okhFICF9QvPMBrD
Tn42ic06uKGSR7ZRwPBaA4NbAQhTYsfHlaeNS3bM/UR13Dj2/TZ4i7Cexw+sZUWK
RHiwVqiJeTZEuxpgDtkTL8GKH7raCMxORrH1pK1wzUkYvbrlnT8bukvj1WIU7pRE
tXtVfmKe2sx63urDsiov2QrMQznjgOrhbImaD2b9KpBaG3pg/g+3vj1Md9bOfKSz
lpQX1TkbOsmML5OEIbzcHAZUot5cFp3fBaG+fSTTIc4eiZ03VA0cOHpSWdnWwOIv
OlkPsdOZAq/uqQPuin4JrWyRfD944xBa24bKNBOTGLn2WE6IawVoFg+AGwb4caCl
24a302EKC9Rp7U5y0PL8raF6NldyVazGDlHcIWMHGzCIwaJ03nWCbUvBQw9ujJfy
yEJZ+svLVo2RoLYiQRWr2HEq2RQ905nLDFJKMA1QYTwjVuXyK/rA+WB7myNWdzw1
c/QJX42qL65Z/GfFQ63Mx+viyZgXMOLfL90ItNmnMo4CsBXUFsgT00eDdEDmNlQ0
VTOFeeRzRXXVFJtowvlKQXUPKwLgYFfOMX2aDiIKDsz7W+fdSuxpAdwhjUTlcGLU
LAywoFimeqQH0NoTI8oZ04JJxbx1XGL2mSfi793m1P8H59YLI2n5ZN2M2Zh07mFa
oZ2KsQH75ejhJOYKuuDHLBM7mrIEypNeCrlsv6eSOqfT0CzP8RBq7lEK8ZavbDcD
lh68WvgrA/b3gqNi74JH5YvQArxP3uG6iv6PPDbUkaWybNmezD2IegqSTaJPY0P3
lMPdj4wQ4amRzzkf/LFUlfMpzzZqFWz2SGcF0hir6AOAM2+p/M46RQGVNumzM3hZ
5yMhwY8j+a8FTVOPF4170FFo2WEPtRb72PNAClC8JEpeoYzP8GuLHN0RZkca/8OS
iDgDgP/i6mP1pWC6NUlM8yPjcHN0vxTSoeCCPnA/Hh0NZjc5ku8tNqubCo6wmRvS
IX+BitodSBq3dLAqirst0OIrQy60jSeGPuF2rWRvHcs5O4IYPp1X+j6XCNwBus7p
0Hq/lRkM10iZx0WgfYqCdYWQQozjy42r16ecIHMTW+XnT2RBCvwBC6Uo1dsRXGtz
2QuhirFKN/aHMoMY2VQZYz7+208DMI5Nod4UaI8AmxudVP+hHKsOyVadqGdEaWFi
gbzHsbDdjZv7R+CwdBu0VtGESr+pSbAmCsqt2O2a/3JN5/LI/HTux9kUoAlEH/bY
27nKkfHmbZkdJtsXQk7hO0nOAN18nZAmbhxZAm/ufROrwpvCkmdpjHebwJnhmjpa
MHLggQaEar7DFQO7f+TOQaNqwxfQ86qNXB8d/rRxW9hzuAtopZIHOsSkHD2K2pxY
5+oq4WK7rrIWRPaLoDHbiCTANSgGZmjpvHXVX892Xrc43uJA+GX2jB9T/GcAyC+U
FVhA7ez5tAavkJxsIFyYei32YI2UCSczf4MRbThNV+cFL4FxxoI1QGu/OvpVTQvD
T5dsbGIdRqD4a+w4WXhrAQ61k3D2jVGL6pL8Dz2pYGMOoudMZkIn95Mwez5kCyUZ
+BRmdA5px1NXPAWaaFRM1VBOjaOrxplyzTeXJRPRBAACIDkzQwrkgic8i8b+USHG
e3TE9hdBEseXkNjdorlKs/GyzyjNRMLYImGNI/C2EHGt7MToXLmA7+Sx0hbUi0pP
tCqQus6/HoXEwZiHjEgy+9Vl+YkSLQy5aPHnFEeWWxoayu8jyxxEedK/v1NFypwn
jysUFZTSAuyniLk22nvofWLJQmqgOARvbUzipYyo3W0pZ7AnGuWUHrpczmhoTkXj
hTB2bpP7mhfHlV4AFlMUDb2wSpa4CC/jy5BIJnz0QxKXYqXCp9H1ZZq1Ls5Dceiq
iGPK8Fn6uPr6qNuqWSh63mhfu/dgsO2ZGdS7iakbey18FLFkSh7w2BZmyv/jRfc2
DFb6mPl7KenzUiWfqtyfUrRYPjdFtMljqsUXx78T0RxwEpmtXCR3X4c0XhZ029g6
JnBBbFkE8d+HsAruLHmhfUK9eaSsM+gJKcdifLxohyk/Kba5Q723mcZL4Q/GQBNy
pHCph19e7TZ9Et8rFhcslBUZhtlWeVmjhTIv9dti3TRsyBYj0O99WlK9+pALZ/Pm
QccUelH82Wzsk8jyJj46YVgEXuqT/fqwdTKM+ctKn5ZZchi1oFayPPD0fFDw0Obg
OybUkh86Vi0bUW7TLnIgivTWeP1GsFLaXkAAtjHGXXY0vXqW56PssepMxJA616lE
0wwIW7JV8yXT/hkLSKvDQ/hoRB0OgZVgM0vzXQgKatfLqb3lpDIbZKjQP9ZjPSFx
Fo3H82cEbD55Zx4uX/7ARXQMsmJcOXaf8VY2AW8epX7eIN7gV8tcy7hYnnR8YPdx
`pragma protect end_protected
