// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:16 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rL3JTNVtiQZ6S2SeZ8rU9YyoXrqPmbQhKWoWOC5WGa81iSM2tXqZydgAlYFzcHU6
NBC0l49q4++6iYSQyx2M2IPtkgHvTMtVyU7g0pLionISh7yCECnGDZKIr2VZ7u+m
jYmdGntX2m29A+pPF5lXkrpWvYCY40DCzF0JmbWta14=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10976)
C4Sr+trjxynJyI3GfpEpicQQodgybQK4f/UB90NjYnr7mgDMJh/9gTenJB1PC8Px
pDq0Y+T6fqnMOzE4n3xh6G+cCuHfDJzqKWmSDezBF+04pkHvJO4SoO+RjhzIWUZx
/H4QcID1FV2DaLrPMkTAOomTwTcVZ8ZmGjV5LhCqM3nDGFh2R2IIjkA+C28YYs6t
KXcHrtYvgjTI9Hb6XepjWlAN0L9aPGxF39Q8hamd2cOiFIq9ru+zB6jLc6Pa+EV3
Q+xq265KicnjYC1tnYsIbyXUwrBXyRbWvMKIt2yPTNc4WcSHfSRGUw9hcABz4DTf
CH4WU2JoIwvd94nQR854WNRH6mWavBiGCg4BPhKUAENaP/gHeCnjzrncRICcU4wX
CotWezdfb4fBhhIMo11QOwcnJPeXBj06muWy/RHnQ6NzQaPfRpI2ZZdw25MN3rfL
FHPfG4CHsfb7WtYbff0s/d+0IuBWXgpj1MZ5biNY3oHLdY+8jgM8Rw98MLTJwzNk
qkXNMJMUXvadwqLx4kI3RC6MJVTaR8bessPSKa+A5IdBj/qYYjsAYigXg79n7NXj
7AfH3Q+lEFraAUzG56Hxu5UowhyFterxfljkYP6b9d5cskcedmOpsJTOPYOH2835
VLy/fw3ilmxX4I9LjQp6aow0WU4g+bv/2PtM1//6T3ScYsX5CtpuuZO0xUxOH9jA
GNcFWhc+Tg33UxelOX0d9AhxG7u7HaJ3YJMw6ExxlCIVgR2ABebiSjRjfEZUDjmo
HuOdfN4NIF8b5BLVwEy5kJD9ZO3f7EYwBGMK5Innf90o7sE0qDOfiJUNMzhweMwQ
Rd5jnGZDkGtCoDTVW3+KlQ+mWBy9z4Aqn/1WPDyL57ZWSNkeqprATExs6BBQTZ0u
33i85PFs53CD+VJTf21UhYNJIdkONScnQvuDE4lIknm+qv6LuvrYhR31mnylVpaL
Em56PPTXG5DNLKjJMtyfEcmZktmsCioIeQ3Z62LRzjj+3cCiUSGPv6tBWbiuxKJk
DxcrcwQMzZPHVME2+Cc62jRub5VFGlhjztaviLbTTsStc6aeK39sWTm7nXLKIlgI
Mpq5lAwtSBkZxHdXYHv3NNsb3B4bzUrp4I95TsCbvt4IQOLUNEpZBJMXPfEp6WwL
r970w/+hWPRa09PLw5V6PwNQlIkZ0Z1Q3PV5oqMPQC4K1YISpPAohdPKlra8WOMs
4OqMByC5hNjwJKcgfp/huUgGtf547TRA3UQTZyuH/pYgmptyFKlMF4pxlOX5kpec
AQMj2gojTiX8xqIzTp8kPmHyu1ZWeO358dYG9tjyE62smN8ZSp0Fjws2Gpwb3UGX
iRTx36JBSP0z339y1O4hqm9+EHmmp/cdVkLuLkYT+O+V0CjgGuoOGY7++A8edudo
Elde9REK1bbGf4oXg6WmjRshh+YLn8mjp/HnxW9IfrcNDDVX5IXNuvCI1TwGQj2L
OmtLNopT1CvBgaKdfcfc9zAnyGr6Wj7+qgKkS2vAsNrQQ/mmXbt2Wp73fmoqJRFz
kAGIEqnoVDqXcjZjOoMVIke0lBnEeeTVt5rrrLR8gx2AN1JWaBIQTDsAAyP8Ta+c
KtdvJ9Fn3WixZT8Mh8+e7TlvDfTag3HEd8B5aRvMWL758if/6U/yGrHHHE1h6E5u
yetoj4Ccw8KWSTTDpQ6wphLynpwXQGzNhCKsIdEir/DOXQEQyxa5OnGetRY2USRW
zZONEb+GSMQPN5bOw9qfHMByArJmfNk8oSquFMAd8mVkRsVle3dwe8w21JiqZT5S
uH/kWVGYN7DEUuUPDCGZzwMJD37tFHL4bn9t9cezo3gURBCXENdDgqMFvxLpQW5J
8nYeISs5fjYPFCB8xh1keWCN43n1qcXs4JmL3z+8gnKgtaEyjr3NLJNJgubd0UZe
eVd9gOK76ZI8cGZ58kyzkRvohSITgDGxcdod/LpmSlJHQiBBtcxIiq6wroGdwauK
jtn/J9MtXYg5pVfbB6sfAzAF9yPC5qgpRcRzdCzhUB/SJIm6oXxOpI0OX1Vj0QYd
8Y/ITg+FacE/ewH5hRTjSq4SMoI4KVvlUNramBhpSlOFhlRO1QRbNAP3rrcfXeAQ
MF08jfN8FdSvLlxfUQKcKnhJUtIuOK+F8yMPE3BBxsaJKkH7XRZrd4GGlK/KgjfT
ED9X9liuScUAdfssnPwRp6BGRemrF54qMkO839Tl7mQW3G7cMPumtPNj4son45E8
3W25XXFwfpN6B4nrFhQzVQOMZ1EdegP/m98AXf11GzSLJMnGfRPaPaww6lnwC65B
vo0mUeZbyHcmqrBhNaqTvOzwkD3oxy7PwNpcolzheEpSAjzpS0ihVxHS0A/GuY3e
CocaLind4fKtsoUW69gR6Nl5WyIOEQj2+7KUOMsRaL3zV9QN9NFYyedapxozWyno
2AUbUClLriz9YwUMdExF+PzUsm6QpWXH/bDrbnj5ol8QPJIX0UNnNGQLMm4b4orV
6bLdGHA7dGH8NjVQBWSVO2gG7xr9+sWfv1raGdoC9ODbkdc5Z3YJwFYSt+sxXVQ0
4Jymxut/5ZzRUjAEvf8fdHCxce5EIQVFP8o3qjoZ3omIhjjg1VPnMCeWB+cgL93e
AlL5kotQAjGAxYGVMcJa/QwhnJcydwqI9kMQW7Mi4RMzoRSnG76i2JEdPvmaXsv1
4/Ad2H+08QE/XZ89O3ZswkrOOeeTQ5vCCjt5J+PuwRrW+r4nz6tEWyjRL5VnQdBI
K5009XS4GiJbtXgspt3Cr9gJWiW1Yg9ezTZK9gj6hhNcwHOoZuuSHMtHTBfzLnFf
lG1ojOn41M9TH5IGOD6L7PhxlaeMZnICSlLyKMZxyqjBy0cEMAdN7u7TLbMuaeqs
LfTOs1r9b9z8dX7/P6rjs/+7FFz6eJZ9u5bO5JuDvxegqK8hzzqzbWRdZ6FjRzYF
2GjrXbj1+v9619/4gPy4HTIqM4FHVCBMqY1kmDxdI2qW6B1mSnVNz6VTUYEpi6z6
0p+Ta1uff+vPe9UbXi3UwEwF5qnRbS+aySNgVCFCVn3hkvhuHoiEbTI3zCX6am89
/NhOOlxNbqy5X/yF0HXNy2U9+fL+zT9w/7bgOMbnAhAQvFt5Fmknia5OaFaBoi6g
YkZyjCD2d125XXo23D/hFdL9eQb+hmKdMooQdwm+WCbHS3EuUX0do7+qm4RBFdVy
+Jwv+8EnH8TL3ZHf+s6d9gq2YxM1uL8qBk1iOTZMK/H7LH76uhLVDO8fUI5nyYxc
vsy7RfLiDqnzV6q6Ds/0rqjobk/+zPQLs5o/42JiI4uNWyILPMqGqIZcqeV8Ig1f
kpr0J8T+osDK499W1l3mGjlQcdcT5yf8YapmJUvncMAuuJ9bzRkQyH1LyOYx9XzA
Cex2S3XfnzvuL9nT9NiInY8tByUbVnTmO4Ti7hKNsq3qzHEdilpHtjA2sRaWA0bv
kkha20CXxgP2I85BBzi4fs7a8PfDPnNAPSa+Krk6g6GfYgRCGC9V3sppmKStsPAL
Gqo4rEPP8mL9emlt4WtgagE4RDFM5ZvKMOPgEm+j6E2gWkogwiaTk4MjhFSpMHUK
RrRwheZrSCi56A5/PQFfi4j90/7JrEAZJNAPX3yZd4/j97f0IYCh/7l20IfHISBd
O8d4oY58gBsakaAJlI5ldfhPjRWL0VkUGjjWHumehWi9E37xC35PdimdF7ZiQZjX
CJhFiUj6WIwLx6evbZY0Asc9XSDLu8UykMEsKiN9GZP5n/vCmJAcne6m8fhYKznb
pagIVm6wPagPWSHY9VFCjDw8vAN1fcoNP2vCks5ExAJcrAouPkqwohp5uA60mD4Q
CV8JhfstAAbcAGUwQeIp6FvsD4FAsdux5Rp1c2BMkeowdE8J0lfHjdIa2qla3Ppm
M4GiKBU1qwaytTKScSmhx1D5NYIQs0eFEINvAk1s6bGhu0jJjDzCj6Na898Oyhwu
R7jPeAJiC8U/EM5Y8OONB7o24fJACFmfKnNN4u/Bc2pPWIpWzXmDccxkfIs34glB
vstdjU3VBIbdz46O8ohfPIunhelaU2C5GmOjcT8c9taitcbBNr7T0O1fv0XPUhkl
BPDnKYJjQ7wsS5VFcSaCVY/XzjwWdw1I8aQXsvCC4D8B7J80W6m4ycFnqHmUbh7o
jgqwmSvEeeHyn1tG0Mrg+fRqkuoCjuEFXBkA/Ge3z6nrDN7upIYLVjO9u1ShklSv
mxPTcCAAsm1EE5Sdkum74yBZgz1vNvhx0YANtI7J6/RThnqnSVjOdNYpQM7A0OFh
oIhtSVitRJMzCyZXmuZ4lctMbO7Fq8gBuDjcLQyoMORVDULo92J6NiaVctL0QVt0
Q3TFCJaHcEiOkAdBn39GNVxpu1nxdg1no/Oko4qMicsZDSngnqT6/SntgYM6eKPr
qylj7jVbHTmrt0Je6soRiXRG+HZqjAVQ0u8UYrTMxMQO/3LS5Ct+p9bnRfNhuL9Z
jcs3vPCJzcDKDC4AfZ9R1l4WSAaDtAiHV/23Qb0YVxLbcvH555xAdcT5MiFpbS29
W1bWPpUEudmXXHy+5kFTcCOY+uqO6xE0w+MkHGAJXongdWIv8ujUI63MaSK+La1Q
LbGv8Ei7f+KLkaDGlLgZNDfThNsvZMPzs3/utJAIS7QPJ7EMBks0gkhHJkoZh5ps
68TQ4Ei5ERpiirCWN18QTq8ydgZngQW1QrsvA0ZorDlSZZz1iRofYYTaSls3JW/T
jyA7bOqK4aqpxh++U6Ia3EfmuYCSB93FjggbAC8fqeJBe8Z0Fc0Uts2JsxFcbZ7x
lj4ZeoDlohnwhNN5NT+UMrlOJOcqaUvRBYUl0ogjx/XlbTE/Meec9Ifr21JlXqFp
hcimOZiVpeKYeueq1g109cXVt7Upxr6c8+Rzm+lsa2hpCu6RDUjXK5LDMpKTGnBq
qRhhOJk4COudLZ66irA+GPcAd8s6xiM+siB7Sx91bwLkgwIHuV1ull6PoButGqcX
dA2vOrQGF2BPewj+6el1a9JiRJixsktr95XGOk/At3DrB6rXCf4ZLzUKYutl08Uy
PM+NPOFF9h2s7qZQhUbb8xBrAT5lOQUhYpKSpE5DYseNBGkt9gxGXarhmuqqrZz7
t0j4Riw7WDg0wtguZXGznNMiXJsgzLNZXobztPiIg132/itTlm/f5Qs6gwdhba8B
luscOFkXW1olS7J+FlHXCsFLBM2BjEira0S+2dBJeBsO6tZH67Bz6MOsXaWsCStP
w5w2UV7wGKRzuipOh5CPQTfYSdLKcCr+cczOeZ1pVS59IKUVGAqFhYBaMkGBqLmV
coArl2faGsCUSIuZksDAS7a23++G/+/Oq/7HM0Z1Fn4qagJEpiHomSp+8HMOYIxu
ziXRagCGKobGsuNn15ihQZDQIfSWiNIeF/DSZpLcfPxXsJtsli5PzhAMJEesVSvZ
hOxsouO06RGfmiK9ee9MIsc/ZloPD2HjKFw9yHUYj48nXRorb5yfgjifNyJ6AAe5
SxJwr/ZCXuq7qbkw8YeGZEB2+gC+H7ciFyVl3G/J8XXhAnhGsxr1/hDsiiHp6dur
GNkoK4HEYAeInVCZcKfuw8xg8mY7Cfea1EOibz7mjs4Vm9UTM0ZHJUCq0sojwf0D
AePC2rOlxOUk/MKr7MIoLHyICMGj2KY4z4cX7vc5c/nXeNrsnoy48ZTmsn5zHo2y
fwI4o+TR7oQtTwbty2iF76hc38XWOuQFTASGJpjgOaXtIAw34On01P5gWTqfJ+28
Cc/YDXPXBPNHXJrMZ6T2Xpkr1oqk+JA2Kti/o2Zb6g6N9dz9dXf8Lovv575v5oy/
htfsriB3AgaBzO2g84XX5Fmm+yX+ScTcP4DQcfnV5UpmhXHmx95YR0XDnV0PYInj
aMBg4dJUi5NNDAXijhlB/vaIp8sTCwAPhQzEvKWro1fRcH9h5BfMl9pUGvBXuAum
WEefa11E56br+HmrozyQaS1OP/1kWsrB0cRjwT9GAjXWc0kvKahBgbgjlPoi3vm3
xMeoTGgIgupvEjaRH/6oichESAcmSvLUwtvRDRInLL8Is4rUmIWQoV+q+NMMZr4T
jyRpAsl0rbxCO0UiFAsq6CdgOqTpM699tPcjSGwPG2DkglgF8RdEUwbnE+KLdS+j
v30+HdFCCNxtY57yt9oeU0tDOr9/5ZSbgJbinrBWEUAevc08o5MpFi5+GZ0wKH0I
X098Y8h8ycqRE/N5vanDaSd3yjcl5PAIeU6c/d3/miKsaSXhSBG07Bx8PfAO2zDX
oL8QKZtbMThWySXEyhNMGZgJjJYRmaANNQEZfpjqMfKVkvrMxBtnkQKvYpN4mS8I
hRmzNkSBDYfAIt+kGwP4uGkiNcNX9bQu2Irirk079N7Vwud7QjKXHK3DsPX5gVkd
cWVzX/yCtmh1RIxTvXgRE0sK9peoNbEnjEMqv8XTrbbMdeUAbP3hzOz4v7ISgFFL
8Ccy+Fv5WuVwwX6RbDrfKKVzb7kXAwtCxkhqaJRdWfyYzjpJTdq0jbRsKeubxFVE
gumZp+hxlgiwscViaxDTN+IEwS1Q47ntgAGgQRbcYNoJbJxgUb5pzDlWn4rjPYoy
zbGDFPhHUTF7pg95ieQqEPv9zNYCEO/rzrWCh166gJzSBDs97oCwPqZjvJ6ecEUk
u4cju65Fj5FzwuW9MtLnGPjM8PhhH5aZMX6f6clUdnWuMmeeXjtFq12hMKo1alzJ
kN6yRr6zqijobIxld+H0szm19ooWI7EIQRBoX1KgDt+x5x4D+ejSaphVTE+gv4R3
a3gRfT59SUILtWCdmgjsxxgqs/lnLbm5Mr4QJOBb5Ids6XWo6yygHhticzv6t7/R
ofJqF5cn7cxfW1LEtiHslLXNMr7Ps2Ptbd9eGju2tj/dWoG7EVuOuS8MO+0aKDM6
CS1x94EYl3M+HeUqNwTG0/Do0t8oTjAKDbBI14VmBueexQyAsxzDsas8vdZXWWtr
G0+kFnKFHgpzZYnUMJ0i4fuT9OyV3rw0cOsNz656GPJpSbzFWoCaCnJtkNd2EQbB
m141YC6ep+CgCap/CfVaysLiY4MuHPZO4krDyBTfaQQ35jmuMBl2uJCaEnkAfvcm
Tn5SzJvcHFtZRx6XgaL2IO5TezpkZPSdal5UFFLZ6rz8blvqbdBwCINET8xn8jIl
+AYdPwwsA30rRx+LN5KeOGjUMeUYvsVzX4dDOj2OgbRcft0ehuIY5rNYUDqYqHWW
LScTiIq8x/RYcKc0dsJ2vtA6p20UKHdbdWIFE54qY6TTbsnQ5eJ9ve9bGnZVQRep
ikKjIxiEuSuP0G+xcNRNcDd1hIOyRfdX5moM4Pr+yZHjo+6GEuntiuAw3v4xWPw7
a8iONVPaILY87bYKcoCHBD4TlX/EDjgWzIW1ind6bhvbV+9Glv5incub3USOM20g
JucXtzEuEnQnzY5bBmTuUUFfzSErrna++QWjLLuWyJ93cv3DxgIGFEB7cLUZWIOA
tXZ/C9DnmKyzK0J1IMe7XA8kswxZO92JE9jUaaoPc7za36moIf11/XK5oIknceoK
Sw5a+sIczoZJlL6Zqi+iogb+uM5dVVyT5br+sWPtmMOBoPgBbnyHv1j0ADdoJz6v
1ms0WKWJJPSzMBMiKz71mqmrQcGf/RflgRsQ0C1HzOfyuuBdQI4T2EVH6afoR08e
CXCuiczNjzAOjQcylVp8dd8E5RYs5w8MP1upMnawua8yY1ZGYd2Aavy/2nyOmK7+
nqOh1CoEMW+zfWrQFX9ClGiQbZMzE+4gaMRU5IyVfq5kJ96/BZvxjJWg5QV1uldu
7VkcOWaHddtS/qi+Jrn8kEqxmIzvVb4dC7QyYAFmsLdiSGfLiiU4pU62TGhPwzlT
fuAhQGknle4+UphtEikW0Zkt6UYTJVUPbtB56a67tqWU2SOZdfP3ITNllHBzUQWb
53N4pWjM3aEct5QPd4rNTz9aPCt2xLi1c3xbjNDDH8DpCCExOZUDla/os1Y4TJ5Z
IZ2+xPaodCUdrmNfZ/LdQA2UbIQWT318nfPCcOFv9jxH6YNrZ2ZW9+U61mx7g1q+
9w97e670JnatfBLRTPptcpL1z93D5E/Qh0ZZg8YlzG/KUv461Jo73R4O7oeP3Uc0
W2KCkumtDbgX5xHlliWKgiba9D/alI+Hid70xRterAwpRkSmZqU87TpLjKtxVMjg
7gCAcaOF1rjsABhzx0d0ob4DNPBIpEXlR+a7/tgoUXSuFzTGV9DrUT57GQ2sOcBd
lM15MeYlsynXOAOe8VvElN0DRkEFT/sozVkTqJzk8JMPDNm1aKQd2MP+urO7G6zD
ZhyBaIIp7nZ+q5OQtOTSy0K/NlFOYYqUJj9CCJLl4mBdSc0xYaMrWatlxN43rb4V
1hFWnWYUwGQUA00COzfIawXCdYBylYO1PaYuUvVNyMBQnRAne0DSJUe7LvpNlFCp
Qv/y8A579fWP88YLqqIOwxceg5PFfjJzoJ63c+pW62iDbyOFbJADl/o4btVs8t3m
9CGGPk+fuVtoWXDey7YCgJ4Xj9VuvKPEjeFQmiV/7YaJAxZ/imYgE9hIs9ZMd4yu
rZXd2fZICeIEn8xtgRn1r45Zoki2ba2EY297k2A9b3V53us4ghYao61v5Vh0dLkj
lGWeVVBk6X5SelqVYsPctdAQJOG/9m/ahy6BeN8YBjM6MDRx55U2JHjAW8qHlj/k
J5iMf1dhewcGYG7dFibL0WwhUBM+Lm7NOmw3CVgrN5vYt+/V1opYlI/dZqQ9H4nZ
FY0mFgkNjwxgqSriJotzz6mjIwgo645wwIQEmr+SnMKq3iooJau9cxU8+ugMkd0T
oLb2L/3mIHNNtv/vMGpt+fEhoJJJVmCwD8JAFbL4kkaMT/FHcvIQFZOmfsbSCIEd
f6Jaqx0YNBQsQEbTsplhW/USrfs+ua9kxFWz7ZnyfD8adBJwyagRH73t1R9Q7GvR
ZnH49BntoQesuBfer+gdNwj8CKRjU9F0pNsyznY1xaDktS1vdG2bDBANR+WfO3hg
hV3FvbAr+PH7RH6CYkf3edLmUvu2L/XJA/GuuPcrnkuTjpgTGOyDzYwoasLjdud0
OJ7ypK40FVQ/00XSh8J6ZYmfFqF48Zg2J/mcBbFfQd0m6NsMdc9bQXBc+FRYE5BM
XeFxBvEMed17zzjlUJjHdok/LhfyyikE2DpFLclLoVG32ZPn5VjeaaMa8yG9+mYt
bNX88xadJ8Sj6XhK5jqbZdVVJqet0FkQLSFF02v3OGWn4Jjus3wRKFKNti61bIHc
iDxd9XHhtoZQcyspE/mgmqGFtagAYpjTxbdh+lmxHo9FntOMlRwORdBSOOgk/2ef
a41bfW6rvrwfAn2zJlBKXfHlKJN/aPKRG/HMdpdz3C3vdlEzrT1aZz0cPiOVvE5v
18Yn8pnbjNIs/ltniHC77w1LLDaVac/hmlMgbiPF0f4FFGQJUWKzpncM12MWZogo
adU30K/0ZziZnQ9NV5l/Rikm/bILBxoStKcOLRk0qXfOto2Nm335gV0Ns2nfIWG0
M4fR77TyecE0MDBFlZFCFGrERUAtTgA/d/n+pn31Kkt8BLNn0Zklh+3XKSJsIjUQ
Y/ZFgSpojcSiZsXDQnl7Ke8FhdlLTlpVNqhaqiPvbLKVTUNCgPx+pJ/A3faUqCLO
kk10+K7KL60Il2VbpDR2ErZ6wN7ai3vHk6RPHldgxoPF01p48F/QvipBJVr9oP0b
Y/VIPm7P/91dqxSc3C79Mj3SU641VX+/HMyTkjpQSSBQYFcdENHiqe5oL/8KUCfP
4G8M09tbSdu+w3pZd1JTWRsGTcxqhECq7Q4MHYAg4+nq1wnCFSn1hIdkCT85KQ9W
y4Cj6B5SLwCa7q4l+8iqgfEojKX7ksamQ9IGfzBJKe4pCDNRN58Sw2LwuYgqFSfR
JANGUPFrQ89A05bnPbc2XJ1gKq6InOYkMehpbkpiDEydcuEmAr6Ebe/0/7afWw8A
FJibhpCrjlUSDS4y5DZsmYnOvBFKCKHdoXU9ofylJtv6vrE8D9OxAsk4TLVp0Q01
XwCOL4hD7NIdU8/ZGnJEOROh/KbQDe7xKC+enQJV/kVARLhhVjRPdcUMbfc6SxsR
Tb6/lGpVianxDIA5F+H4EoP0nnLLeXOmTizF/nOs9ast5WSnuEetwaG3ICoCMOaG
3eIOeu0Q/KCMQVKQF5rAzxdBdK5Sy7YNnf8046Z8XTqNtBgn0PEKEMCzvPEU3nml
QixPrpfzLB62WSbBGJs472C9LIDvCLO0exCLBBEM/NPbHTkYihPmlmQHLLEPCL0w
DsYUJk338Or/YG9suAnh4eRsDPoSU+rEMxaX+O72ExLpW67wp9TKXUu0cErAY75k
3mW6rZLXZsk+lFkTSzwWYc71T9ZKDT78XI38UBtBekGoifkyvv00Y7faiLH+fnA6
2IsDlufLXHcPPLhGa7i22lPEhm4WleqmFEiaD81U4+jjqIqMg3VCSPl9yhxkaP6g
LdmB81i6SA0lrin4YlXs2c81EGSxURf5YolbO8QOhza8BNwA/tcGtoFCzHpK+y9K
AB/4JRlI1XEktTf1zGnEP0sg/ERGOuQK9CePlhKdaRJ0fF5Ui8nd4dceBmOqM7eu
97acdoYvgbKnUjk8g4tP7vYgr0844PwVm7NTC+EDr1xyP3USRNToYf4GCVrN0Zjg
oJFpqqH68QFJF5fvXB4vqBUTDbsJwgeiaZucqeBqTeThny9KsyIBdE/NJUIpk+35
ElScVtmVPeujrlMsIc2fFTn5wp+7EIn8OU+NCVEaHFnZB7KdZoo1FIWzKBvHKe9m
3mRPpoQ3FOOGH0rbk7g60k7cRpFi3OR7g6QZCFSaoCqHe8okg0ac3RWnohM2c0qe
xTedl+alxSGGB5AXVzKomkvcML4Uv1UBv1U5yc6ClcGAu0Z3DyyEwYlV3sM5XIvZ
TGxMgs+715dqy2qQGkBvSGEIJiKHb7K218SWM22lvvXzYpxxSGzupFRTuuKfhN1u
bDkuclGV0vFYt4A9WtFc1sd42SeVpadVhzM4IaQNtT5JFjpszGycElI5Azgzdngc
s/V6MQm3QxbPaRRsBGy/NL8qo3PNEoCCoQhT9ws1SRIEn1xWcwnQp/ORE7iy/tUa
xLRXtKoeE0c60qyWk9LroxzLkOif8CLqAhwDNdS9ovk83iZ4hGhALQUuPHae3XMO
cMfhOSd7RDlVI7Nu7RczEbnoRHs9g1ZHBzZ5CtpqX+jmlitapol00zBIdi1omJPU
JeHyhZXZr9Q6XFm0792Y3jTQf83ihYzHMQ6XC272niAXxX9MOIcVNWUWLlm9yeh4
R0TBA8PnFDsrxZIUDTx6PzMK1nGHAyOtCkqhtL4KNrkzSdkDMQ1nfmuqS6ZvOxNC
NbKmblT5YtCMGCCLUFCTiRN+Wjg5NnlnzQFFt5mo59De+SCRcGdOJRKuc9xROuGf
rwL7jZTDb0PnUPu7X4+LBKC9Pd63MgVV0XH2z/xXRfBQ6j1UXStDuBD40xp2wVaR
pAunyNVro1HTRNBmtrGMqK7USGFogfv+EOq1MFA89C/HoLQ8rRNSW3VIB2F/CtKf
6b+0uJSE6tVuVqgpJQ2w+kqM59nuepSoHmDUAu3K7U40pvR6DD/WcEObIqQWWjlw
NPNJ16dpgYlHHOg6VKu9b24T+03eOAtr/KasvmbJFkW27Orwl7lz5uCZK/R9MG8n
o+VfGU28wQIVhbe7+tf87sTZvCgYUzhRj8TuGUbz5ADLwIZfb6D/jby58DE0oKxL
KMOucaLYna+zYoeN8tXxNVRx1EgQmFMBfN1v6yJ31z3Cjdh+1o8ifVs5yedyakdq
+g5jLR4BcAW6Ow7TtS1+R5BdTIn+jlcHxAMc07dvJSneYok4aTnSaA+3VhnONmWd
VmRu/i/ImmsFNL3AXa+iBzufAfCshP7L+m0pmG+MRJIaIsEjCncA3BToeA2Qaw+D
5rGxWR+kVusocxX1C3QAQUXHllE0zEpqBSkQIkiIE5pdawaxAQKvYhWRyT3nfcHl
nT/bJxeugPpJ7f3Jvu0sqxJKaSPAG9aLUgXuh/5IBckJW5dzMwHcxvgAkWBJBbvJ
c9WefJaxIwNako83NgakRuwxupKDr4xl8mxSjXpLCmXtuVYLTd30gzuuXWRZ51bP
oArXkgZLzn5bhodJoSAt666N937BQN5J3mUvdEJ2rg/pK8Qf745vR4vHgI5bPSOd
pft71ifQiiJgbemrvp+77W9zn5tYtN+/Pbmj72Qxv8L2nkjgNoVw3+V4BCP6t2P5
bF/fyoY308iqz8wH3HKeipdwNUiTzOxyN/nIo1ezc3MmI2TAkb6a8w9chu1sHr2M
aNeKYsEoMRuucV6hlu9WWcOCXbGkbge9EVFQhsc+A/lOmUjrGSe8VBECo4rDV4Yy
rWJWKcT3+nwUDQHaY4vxu+0AVK+0D66FPI1FbNljekmQi6/OG6rnoUaHDGsY23Wv
TGXMOA1KSTE9mQEZOerwc9PPnl/6h+jwjjp7xi8W9r4aIqb1RS79OVh5u1mrgaXQ
BjM3uhLxIfm4lBXHEU/GMyBKpyVuk/9Y1fUzuXMYrI0NY+W+gO9XM0CfsHHpiEjk
+MaXPOiA/tADIcGOeU46Eu11zLEa662Zz2mLWoIu6fVu60W4PPrRsPwk6tmY3tjC
SD+0AoHQCjhqspF4q733QDti8VNmIAkKw4kP/DA2/wxPC++j9M5Dyc/9Q3HtXHIR
7QqEcyiWwntacdiSXz/7KDs7D81Y7rl0JBeWsz+slDGsNEnoJshqik8FP1tP155y
r7fCpnbr2GoEdHEPv1RKKffQtYfWp6DSUPFrEetwQg7GTTPYXcsW+wzKrqE10MIO
+rNs+42yV7dfh/dpj7UWHwsXkgjXnQ0Zin5yCoIgEPuApF23SZhGocZDRH+Vk48h
q7Oeq/dA+7ZMoIXkPU0DELIzj/DPXjvlc/xW0/r/UBRIUEqVb7G5U/QTstzY7e/z
U1HdD1YSGcCxMTRFfUE5ANow23z9siXH7MiTUByDC9qRsgX6FXEBWc3yNeg51yHb
So3KO4bixa5jp3PPVO7fV3ISKfqyEXOPzAE7z7PZKTpU6Xixfg6qcaw0tjpc6/+T
kZh2heT3Qz+dYiWXhK0HCiSGNbzwVdUSpLf+eiBV9XOYYCu8QI3fDpkWGRitOuG9
4Ir8C+Ke9uRfLmqlAbipGTI+HZxP9XPoO/Ny1MvMUQCxJX+pRZav3/Zr5rkopxDX
lTqocIt4PBye/0NFPlhvJ8soncko2UpfB8OCurkK4JKvN0GwEoBMosSfGD5V6ATZ
MzlYRfMqBJQDS96Vc+JeIgCKCo933VmE4pnbXv4cMZzuybpuu/PXPy+c+EauuMXe
O/SaZL5nu/fNPMJi6zLjgT1O2TnXtXS9aaIml+z7dbjC3FhZM2RYxNE+BO8aUoo8
SNwYFr6KZoXdjnwREuX6A9HbejGp2+sosZkRvrdM1cftuWLAw0xu8vctFClH7+im
e3GHg1sMV8ix4X7ofdnExvVNu3FX3Oyp8dinQJhvoYsLMLX22OH9/dFXyKJOrKz2
0xZ1PmfkrCjCWxEHRq45EPg0lNYLe5MNEYspaEmSTanK2mz9sN4whbg0U3EC7Yv5
sNLjJB0SJvGxleQh0bOAil3pEHDrLIWmj0Bo9Y+dMdYxE4GI1ScYTeSltyn/TTPC
gGz+UIo5gHf1usLD65/E0/+HkWhTQXyz3kF+zuxsB93a8XTPfrM2rkfOpJnnwcG1
sjTkP3bPz1RflUa0XhU1cKpvwqbEMpEbuxzA94BMrExjBYmv517WV84434B7ZVmc
/D8vlOXBcsGSOWs7g+8ct7iwpZiDbhEOs2Z7mYEV0NOBzVSUlEZprM75rzX31d53
PEmYAJNPvuP/L1t/vbB+kvhgVnALAlOccwRxZ14ylbCrs/dFbl2IxTg7afmF+Ahv
hi3hIOxK+Fsd/bHCUIoyOVMolbfrhxJHllL49HuGXex5f2N/nwlzjg+KTckbcle9
iU3UARBXIEL3EEUsk77lFZuBprCZnsx0P1TeWlfx/U+L38R54+126XTMfP7d2Wbx
6MBtD9dlPUDqQ7N3SI/qXUVYs2Epg/FVPX4staaFOIVUPEs5vqMzMFPWmiYxOOYh
O8iNaTm2Z69vzX2okSbANv13NE2CyeRNq+iPV5vidt1iVz/CQqCqheSuB4GSzo+/
QAXT2Ci+I6SzSS4w4cEpWd4FQE0K9a8m5zEAR8khXzPWgBaOp102MjgWWYafvZ3T
gT4Bd571w3L9X4ozB2ApyBcXhwikoxnSXBsz1wjGt0mvoQlK8oOfS26bzxf3pcCR
kXpxwe4CDkNQDD241U57iiai8QgXGnjFzIEofyaCZy7JtFW5fzCUEiuSfUYFZKlv
48zbzrhnCukKePx1P8TrDYIGdWYSEc3yN6o9zK5CzkmarSKdHqzXwVWiiDBdW/+Y
+Bc3NOaQrf50163m/VurR/rds70Gn682RbQcLIKJEmbGyVrtprmACzVtQr6XGAnN
WOk6MTntfyrIruA4FI59d6o4JuZmqnNGFv3PWe1beV90kOJpfChEtxFL1vJGdewG
BsTkkyBNDcXG9oCZuWGL1SRLIjPGNm33ZlNzoyfAwdM=
`pragma protect end_protected
