// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:27 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OqS7yMNARfHoVmiW6QHKnCfFVkbVYCy3vIdug+APHTZvxih/8E18OTNIlYsk3BIz
6LGD7fxbNdKduob3UtESjK7HDPBgn1dYRqAZW8sGBY6h3c4XGB1NBuWJbYWLMRZp
mEHJHFukvmZ2/vfuD0lOlwH/RFTKNjr3OziV0S3SDZw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8320)
J3KJIGZb0ZTcNJnQiqaFzfHTZL7s4NkUe9+uzcz+8YHEqkTplHqVRyGUzxBRlHxq
Zf9wkiK2YZwp/fsxD3X5fUBjQSdiljRpSDEgvdKtkkGQLZD6ukMf0sq8h4yMUqm/
uNhD15E0Z0SDmZCtAaMQ5/jsxSoqGzejaY+pO/DFdsdvgVTOtDOdrKogLjBWz5o1
Q9doKKIrhtgu6BmgUC3cMrqe9BQHaraQmRAjd/YXNIwtnQhNel9hmABK7bbf7t/e
Vnl4xtz1/YsRjwpUF+Q2iP9UTL4+Oi3lgPCdDpyCkpNmh85yDzqf60ffWLtnJttz
YNuu1MAzWhzP2Tvc2bfWp2fCgEaGncuyuAJ0FL7OXTLcjYfVNhvgf92dW8oirzHF
os41l5QbZPqIg3ZpX1ERKxoXGfHfWcC6DDaDulR5j8YIsv1JS9KiO3X7MYsp9wtk
z1THe/9zhnEWatXDd9bPacMKOFVhbk3hyKruQaEeuss/TKVloe7YQU5dAk2BR/1V
cHcIdtOo1ek0Xt621ivVk97jboiqfU0UY8TR46YW8iYvd9Ut/LwD4AIrxPUAEfRx
mdTuNRgUp+3yuIttxC57UUnwlShn96co49ieV5I8yxn2krK47xeoq9gGqNJbiEgD
SNl6mNo4pJHeOMjWHpigi92T9XTj43RdWBczCNwwLSPsZ/ooKQEDQ3mummtwB83g
QMWlFtGcYfRjWYdTvGH63iwZjQ+HOCMkfnQDmDad8H6IDJf9tkgY9Tjd81LVqHI9
+zc3Rozke1hw0BQuBwOJ2J4xVTJHvbzqvsEb5kiZVDmXfcfHMXLBZMN90p1Vaulr
8oftn783ug7aiu3vz91cuVn2P06Yf1L6CttIPox6v43dVg+RehI/vZe1s0oVNIbY
d5yJwB7niZT+QS0YvGITdyv4Z+H6XvZO6CH/NyYzJFaWWQwwwcIbloTjjUTfN85X
Ejvlcz2kgJS0SopzvxKBY3slCwTIqB0roPQAvOzXPLObxM8o6GDsO0LcFK4SDWhY
Zh8f5b0g+0ZpyV2XgIYTdTWV5hGuJ4JQcNLkdg4ub5fx7YcjZ8dInmZKHEFHlmLK
OZJSA9HPj1fP45gll+sQXucckTIS5mOln4mDaT/pjEFnaXqbaZ2bYpsNQXna9gVm
0s4zv9q346i0o+GmNh1kYXLz+QmShPKzOOazksnLwPLXKL/+rVbjbttKax0EzteR
OQkBntvzfatB3TyQk0yDPJJioyZ6BQEYGZjrUFl4J6W9MeWQPe1VvM2Nkj2N7TLr
FBUu/dF4vr/GTKSUhkpJY3KaLwaHxG3NMhVA8eSrHwY2FwF4zbYBWCd0v25EWZkV
IoEXMe48q4QXINrsgXyM3D9cicnfP7UTNrIdO5BX6qF0YoePgqo8L/kcfuhgzs9Z
lZSlmbZFhl3jeJ3Qjdm/eylmXSXtcpWIeNHynbtcu4bH5KX3jg5zXjwTov1ZZHI6
AwsA1m5CG19wGIE23f7Kw8n9H/6c+f8B4pnGL2zGVypqDnktuCEQxX5wolaoPf2H
GHl+owEAa8OWkWOd75aouvWH2nHwx7FjyvE/ZQnlp3ymluiyhVSCvuDImts9HzkT
blc21UC+Blk5hvXQ7s+QyFCXOShYyIZv8Gk2kQRNKmWz1WIJGv8sOf4AViPu/pg/
SktrT5/CMRN5DHJV129uNdDotLKkRpCHUV/SVvIG6rl7OzLQAdJFsHvF/bTQjLvp
rRlqOsLBVfpAG6k90tkrKHom6dTrDcdftJYEiwn/nCibRoOalSgLr1bJf6MxLyFg
E5dfG+mf2/s+EFZbVUe1MEQYgQo/GTg5CK2+2Xo2m1ul/wprlp0MeMxrtkMEOb5i
auUMLPuihVChoxq+71daoqRXyZVl7l4gVJ+ufLb5haBed8urx/AzjyaYADq3IqF/
po8xcf6mDPYe4O0vumETDog9/VGKxAUPVCJFTzPIxEV1sGgL8Ye5F/dZEy0qQsP3
D4JdDS8rfnZ2dwNiqKk6MLwuehSFp/I077PnwTpgv1Jpjr7Aie+X7pgWhtPHu3J7
h4dOXk6Pm+nSayjnMUWE2JRIbYYMlHtKFX5rLVwxQP1jYc0c9e4mxsZA2Z0nGX4J
kfqnlnoOJRlxawm8d2bufZYM08r9yJeJwwcPjCjSrH22ag9nPElPmc9xphql7+PB
u4yZxI4YBciiOtOhhyP/aZsmCdFb2sLvRlDF7tq0LgfqseY1us8tBHsl1bWap7L6
jnKaWcObhOOENdYX5snPSGEAHCNn19AdUI854j5M0wisIVpjREtExTvPjNXAWWGJ
XOEFg9Neb+1CthLzhFAjvP2ZvZPz4FDWM2cCxkGIk5s98Lx4ce5A2KpO8tzafSOu
F7Vm4C3DwK18dCM6HTU7Hk1fFtn6di2siKHPLh3yJWzOzqpEiaPCFKsUBcJEyqgE
b4SFJAjCmmyVR5pibr/26oLALDttXfRVHd71BeEemnvxr/TL4AxD4FA4QNS4KlU7
heHAmXoVcFdJM0ln4/eIP8eNfivCwOFkA3BHZvd5abo555MSE8m+aqHPePOP5yXr
9W/ippHOZ3xy79STHFfWI6c7zcANM3arbH9qqW8Oz/6FExyoGCbZtTwdvWEHuxg0
65gfaA/S0+HIyq78Z5O7iu266DmoN1gJeFlp5BOw0rgiMfd1vmdTs1mt3illWCkl
cxadnHqa4jIRTeulsZTHwuxSSOoMJ/rBz05dFqMRjOiN7Nq081NE4QyezKdmKwsA
qtGk7z1Q9kvo6qUqY+K97F0tqMcGLLkomv962MuLq33WmBSyBu3cabB+JasL/NwK
ie3r3kaMp4enQL/2lSw5BM9WClFRpNcQCpOG5PrEsCIEHmDFci5rJSOEAFlZ/shR
zKbCljzy683QzXCYxtAmFBEoZuLca4jSovDBXPne6r/qvhuRaOE8sHLjUStm1NKx
DTqERDQ3iVuf5Tisf7zFDKGaDDCKi56HINu48w4OLTdQ2KMdOxVxK0XMm82hDhBq
77ISuy9IhjD0h0Rb5sZ3PRQUu7W6I7/1B4FjIADD9vT+1C45XtXhz6BAW5iQoAot
HmvKd6h7MvaCA/wauvDXpY346g4DQP/rFBmSgJ93zfwrNGC7SNwFGHT9gip1Axf4
kf+63d6krzHImKM3fUpAhgsPAUTtWfBeEITv/JaiiUs2j3B0DPTJfqaqYqGNkDgW
E11O+XgAnpMz57sqNvyFBb3aFdfXx+llAxuotaYe7922qvvWjyCSzWTYpOMrI3My
J8t+3ATYGmM1XyG1+txOFWPtGB9AT+uTxbtTaPIO6xksCdNGdhfjsFAZY6lKYQlz
KDle6lwEuRfK86lTwoJqVE5e1w8irxiVrcbTtP+bve0Ta1n+qszmLIzYtReWf4Ni
uDvTwJIEkr+EuPnSayk4YBhHcCY2e/9XUkgvjvB0p6kc+lvd/bc2MRdBoICZQg1y
jXrAMPNn01PZj63YKkEQPdgsdAjgxfBgN/xIS4RZq0chHo74y7Ewb0WNqhS8WjCA
Rpp//IhGu2FYb+9DKsHN92dN+Jl3Pa4+JbK9uzJ+0nsNEEOLukZDViBfvBFEKmWs
bEalU3M5riODhz4fOXc32WkowfGsstMeIhfP4uSJJly1ts+BD/2qQjB/+IktUWQT
Hehu49tyq4G5hqg4raqoNErflmrGBE8ijxE7MuiZOtHeSlYBrFS2pq7UXmxTft1r
6kr67bILL9S9TrbLRjmy6H5jjtB4JEgJ/4zmH7GqctTpjULX6eaSCnLOPbx+T5wl
GKJsaAMpcaYJGmHHwy2kwWsfuGqMfaB9pENwFpCJDrm1UM4e9jzlWoD3HE6oSJ05
XwiQnecswi91WO7VjsJPkbG5LN7WoIQAUVa2AWovLUYSrEmBDHhZISyU2UaUICYs
kVe88nPquHDWr6huUZ5dUfFiSjLNh7jNLvwHiY+DWWoia4O++mAHD6F6acRU9L2+
mmC89NqpwcVll3XRC4ITABXiXULuNET9qPhr2LPoKInAN6HhchkhTbcOUaQl206y
0X/Wqyft30lVMdNqc02EJ0oX1se7B3DMfTr51p7MyHNyMDM+cy3WK7Wzsz+9V+UP
cDr/20LYc7UNwb7L2PNytSq6iaE8MhLNQ/FHVDbMtZz2O0Tx8NUP8AWExG2SwlsL
Y1fgOpesJjQWGiOaQQpWson2nJrCzK1pj0K0v0QM5hmliVJHHldfCpREyh/1SCc0
XqH/EJX6uefO4GZTP9R4tl9BEuk/EadpGmjQ4MH/6O6axe4VyymdGgNPLf2i3jov
MEFyF3ochh7cg7vqZdErllIj7kG6mDrlujiNxc2mScabdr/XtBcQS/vxmjzBDS8d
u5MFODgIBvJ6Itt9o7vfw+o3+Dv0JuHUsgf6vB/g5JrAnBHSZMejpq8NdeVhAMVX
vxfRpro/dXa6q4YohzpiObbPI5d8sUCtt3HBBnBT4QW77pBNwq5wGOTD31pXBYAr
HOwz7WKXh0+3wck0Y9GopnK9B71rxUoSwDjdul0wjf21W/9QtRjAhGCjq8auD8dq
ZfJQt6fPk+yQXTP2e4Vnw0wSxsx5F3Px6l3pfs9ABSXyG6qhwfEymSFLbchO9OEo
lt+jnq6A0w5IqCqg0QlifySreGuSX2RqsuMadjpWNOMW7Ib6JERsKvvFnbiISmJh
lvqmPmGBSZs6bngnVgpNVKXtMrK/ziEJmNEj/kvnlqxTCHVIxdmyGlT960YNGZA1
7j+d1oBzPM/4+CzHy44Wz0DbB2d2ZNqvJWJ8YBzgAwtONqtNUN+UiVEcsSVhEyww
xCrfQpvVgRZ3rM7MP/IZKHsPpunDv+QHLPZFMbAVVXZ2pgnZHzVI6CHKunLxoup2
9enNMIo79Vu3Hx4k2lHDepNUsPHS3LTUSkqStQGf43g3idnlfEyRNMZMCognS4fa
+9wsxdwzbzCx1h3rrqF0lN8rnLHTSd5ZwZGCjHOidabWCueMrjvmwgXKb5vvRjUJ
FLECtbNhc5eJKdHIdHiYYLgkSA31RZ2cSyoC8xWbs8pwlQkzQQ2U2rkOssyEK2kS
9lhEO8ZUaqUrFSz15gsMEMls1Hv7E7sXzwUB4q17gH2LkeYS5SaBqijiar221DRn
sIKgmPjTZVebZrph5GJjcIJXMc5QX/B80Jzpq0Gmq+GnHB0Ao5UET17wQZdMeAFb
95Sf8HW9Bp085VFMUqeDo6nlcsgn/tQWjMzxL476Sk6BGysDFpAleI5XTvKzbOat
4lSLyQqPRtJbBfERP9R52FVz4zJdZre4SXJgbSkZGLca2x0h3AqPLqgjrXCIWbnr
dLQbxZW48UH2csBLsL+eycH9iNNTJ7jMBxWZU2EHFlAQdtHG9A1I062kC3i++seM
+nRg3ru1/ZJ+ETYzDq/yM7lToTx4dkYtEGXnckyZoz0eRmITDemkFdBNINsqa0Ts
3FtwUGMQO4FEZybPslc52a08R9jqX9kkOBHYV4a3vqVTlrZJgTWN8f9SF9vNhKII
I/ohsc/7BCW/q1VhLsUknoph88VBTkHwKylSxRRT58slpEftVYZA13VJs7k7JPL3
JPGB870Is4Ye0kuNAwY6ABYzezzf3beYE/xsNXo6KRm5BYJ2O0NcEOq+8dTU4tMt
wFJ6hKsbPnk4c65Kml1+wUsn0txwvwYLd+Lk/Zkb/UHPAaTBdEg45YiTIqwPpzI2
+/uvT36daaPswvGa8Kc/jutcGaSW1HG01olW/F1eJ5kXDjs6m+9DVVsfjKDoAiwX
LT2Sxg8s/pcSGaLjpTwblXH+QPaUyEkf7XxzKOb6lEihxXwxMwb52794YyOAHUDP
QTyKUhWJ7sYx9sFbf8vxe6LsP5njhe5oSeChsBjkjES5kaMbH8EKcjz6u24x8Tj9
wIqw84OgrG6SWbmW93na6AwvL8jRpEhLtj0bbTrpk8/wmnpDCx3an1ctc5m+R5Hq
8vn6AMBOg2klWdnCYmQjABWIQCozVwujklpJNK+qgGLb7d1Gy+z+IwrnIclMtnJC
HLouqiVDnOEzoqI5EdHatECyIuUvFcMlvUJW8Vjgy3HZrFDUin4riJVbVOPQNeXR
/TQrAYRcJAj8Dflw5rcoHc/NTDoUcMjvKDx1sachztBIfMwrxdjbwo+yrWKPYYyH
rK51Y0oryDVg/N1jGS8wQTOMcTauQ4VsRGbPg6qAlAL1RUQjZTmAkH97q5ZSxmwu
A1Vsj2u8u6Z5vDisQ8b6k+9I1+2sOdDDYYM4TaeGjHJ/3j83ZzNd+pwdHsJDKMzN
ckCbKOOthlrRV+NEgiXkMf+1pH7RSgBopmbZx697Dacx+uJoxXFrVfFwHb/3K+st
k5WVcMpVon2wIJXuDvVeJ4x6pfjS1W1Gnbwk1IXCZ/novH14pYO622e5GNZDA5eZ
TC7KSugRkr01XZq9Iv5adUdVXKh503nYI1zXqNlC+//mK7FWz/FEs/lsiK5/irZB
i1yAzlY0/wCQ73+s9lWfhs8OHZk56BISQBwsEK2Qst1cDuAO7hsScpkJtzu0dgO5
DECcpZ2Fc8PAZlgz7OtFgtWrfmM5sLAelpGI1LYF1k7JKbw5FS5epHuU1RihamAS
Jhja1WfI1gRGfSSuMRcxygjo2NpCEjx7dY1ARjBsV8K8ediK44zJG8sj+Kg0xquq
7xeLRWTYstF51UHHPpoemXllODa1U7OyQPwuh9PT8OX3A/YTnJT2YE6TgCLWh9BI
gsPK371BfXGK7fCJvgaHOZVCoZFqihFD4dakZmqAR0Tk8X9LTotze1FWjLe7y8MB
C4NvPsnhLLxVT77IZojgyXrW/0x/bNcPmA6CgAedK9wc9ZhXXNagUKiVU+fRTtQh
BsN03n3BMB2vAsDnMqsWRnOJT3SzBiN4Uc2xgdU7WUtMuuAyevY0lq4Sp8up5NXB
IdUOWSMq0gXAjQGiVEaR/js7sN24e/EnCm7NaYEDPVSmAzQPrWOBnzsJOvueYaOi
ZKnZ/WRZQSrWakTNYpsOzD3sl/CxAVxFzUfWvNgSkSPKDDbNpOfI15tNNkiQFACQ
PkWnNrsl504QFEkU9QbHUivRl4Ym0udw3EFw7sHCBRscTEynDBelpF6Lq6FKDS6c
Dq3NUk3jC2ZA3m7k9Z1pCOgOo/aOWiLMQMkNqlap/0woF+vPfDzrDMmqYB2nSUSx
ovUTGyoWhvYw73fo+c65id97j4ADTKlxRox//eS9twrpfzXKuL52SbXwZuxERt6g
J7A311WrJ501oXw7olIWXQ9ihsvoHHWdNfF98An1snMoe19SobRkr6WDvzOCPtXf
nHC6qUgeSEWR/MCXBoFQkvEo0JCh9AIGBezeCK6EJJKG9nAJ7/VdZLT4S/VMteCk
B8/C8+c83vOh9+YMK/RUBJu5TNY/zmGpZHkRsXK50ewZkrs816zzUs0NKZ7LA2t7
T6pGNucjLTv0EwYRj/8fol/QZ+x+ym8r6Jd4L3AHwxf9tZz9Tcrk5Gz9r8s9Jogv
KuAOGqzrTWU/VZ5fyAryAUnFsou+qP+KFfP2FJesyV55i39EMvc18S5M73fQlKt2
McKqn61gVo4+5t3AuRLDGgFCiR2NEGo1ixRCwKQN+HWZllTwpF7gla9YMHyK6BQq
QtkR3bwv9OTzhosPaxrqlDqXZCpPKieBqwCfhiwOMNuReoEfX0Gzx8GshlfF3jJz
M2b5C65yrMJvKdDDZURRHkFZ5Y6s0rhIWG7/0IRaHfrsIELERkmCtrdH4wFTzBpZ
LEuXA2OJR7u7+AkIWE0dOYq9mjSor+cKb5fV5dw1BrtSmGEQnPtM3tT/KCfOlO0c
CSvS5PEoZK5m9OGUfzxL89tE/D861GftolT/BBRANUiilsAJDxL3p7OcfIn1bQkQ
pS7vrIy/81kJyR35drhAtVppakSiLC6cVbn9W+kmxt/sKM5zs4HtQjwdvWs3Uvuc
hKh15tqS74DwCXrgvAVJv6luBz9oN9i/ZsLpgRdvqQm+dCdKTMlGkVDkYZCe1UN/
xWI+DDCD0Axb63LAczoXPDWoWBmN0KBY5g8Dlip+O4Xk7z4Y8CCwk7w5QPnO8ecw
TRsuif3xslR5lvAhWgEuVG1uaXqLrvtKkrGkRhS0PL1aXPdLPRp+2nSH5WCHL5d2
ky7jhkX+MBXtnaeqc0XvxH7cwrEhOIjUXZQWpkK/Bd9zdmbYdLHH3lj4X/guAH06
Pwg7/+a26F9TSz4oKot4OAnFCtcUqBpuUdCoNz4muMqQ+cCnpmxO7RdPvp01degS
l6CY242R8X2Izxp102E70FzHsTbgjKoo+Je2IFwDgH7Q0U5XbgEC+flGZlnKsIXx
UQAbBh1B+nLGg2XqU2FlsZPoboIpvTU4Wh+pNX71GBBBabm8tXa15LNu+6sK0iPJ
uZF803T2qkKlp1bpWYCD99DpzkjOOaSEWTuyzu575tFCJehYskSGjDy1/ZE4oz2T
Jrt1GRek1iWjFofcmJYAOdjjdnGHSsHsilg+P+bsifPtExkbyTeZOto671EgXIRy
KiLvIBv8l9XSwQwKgFkQwP8RaQ5+BINFzRgGq6P1kng3mCShcergXtwj/bC66dTd
LPlglV4apWtQ6WPJXTyaiALYsmHFL4zQOyuVBU+ttaHAs6k+avLIf6UctmWzz9Ic
80E+lmZtFL0vx2vbuv7y3CaLXqUJNQcUIotQfKMKf1vOaWhmD7cGGK9uRkq5mzXh
6+pGojfJimrsrNVDAS4GV7fGmfuQii4iFaNI6frBdDhoUWS/WwhcXIQWydl/GlGD
JCtGRQmHBVXExe7+R+PCjdrVtsebskoxGnxeBKv7xwSQBQDp8hmQVBDTeHIKC82O
npMdh0yz9hqGrzZj1YYdqIW6s0W3NxmuUYpslRVQ3OYOKMAGHG5hsq9RS4WIgcAg
pzrr8kPo+hCxKY6JuxRueHPLlT2t0SFGkf3B3v/IquhTBMxOzHXqqzgbrHJzJ5d2
46jeqfBDaWChTNjPoBBSrUusIGiqgnPIY0Fp0cwluNNbfnqWxB1RI+/8vIHazq4p
/a9v8nc0OCPDxQq9sFU6bg4QI2Nt07IH+bKMyEPqCHIc4swG+NO5lpOgoSzPmcUD
3TbDQQ+ppp50zCtRHhp09KN3xndVTsL8nse+69xTlXQPFfRhzljP5rOTWF/JZJOA
zei7YC8uR/zGn6jzRqzuwhJkREPQbYxtRkPmw0CliPXkPe4IU3+9xqaaEoNidSeG
UN5LogSL8DEyfEmtM0PNk9NeqTUidkMqLKl30WRwiP/CyvW556yzfnKmb94dQraU
/+tP2TwCM2sGVSc1hq62FwcS+ynYgeesnzIwbkiu+YuqWWw1UYB5dEoevU+5q+DR
0hggQH1ckkb9bvyG5IaSqGb66eXK9XcNcFWmUfLQgd9zYg9RTv9/GRjnjhuGrMJy
afr69LwMju78goPuxIJzlXbElISPFI2YfArW2K06yLAC1z0YAZDwVJAQLoTWCdLs
GRYoF3d00GInYwR+YBXX1TlGsDSF6pvY8fYen2R/7yreBm/IBvM+5dKzRjzccywG
IoVHr3BsvvYxY7RCvUoYTzwuCJc3rBkDVuUDfUS96zaxD+wpZJBcEI9dntJUsRv+
ye1gavm5E7dwaaAx3a/H+IqhxCvlaFl85Wqdgd7wor7ch07HCn0gYSPlsSw0r5/r
tGxlDMwGqzRtuGYP30TXfiERCrsxMm6u9O2GnYej2UcRg3XkEmRYix/+zKqvgYZh
pHPk+drKhdQs6ESMjLFUuvYmEos6WPcNDG5LNPlox/4VFdFZIqjDiTGbxeWniSgk
DEWgC5/CWi9TCbVE4nBbZlhVwlqnOiHpFr7vsP9pGfziXU4tHiDYzq9uJRlGXRRu
LOBPDfBvdAluFbZH1n88x1CTGBD2qA+/dOHb8aHxGrPf4HW8khCQJzg0Jr8e42uu
Ko+qhxIiDBOFWbvKbpM+I6y6XLta0PIo6ghBw6dsSSQhD8Mw9IHct7vT0/AGvsg8
H1ow1QNJvFSzRx3kFIvah5aiyQUlXedtxvpwNo5ssKL0tSL93Bf5QHkIXVrwd5Oh
LEvCcG8oYoVBdf6LotEO980gjglLBtRvPrgaeCySt/3w9cmPWbp0nfQYiG5CfUnP
TR8FY9T3TZtSdbyMhZEeZxatgNMfTnJLekkxaPtnp1hUXqVSmnXvx0pv4COibt+C
wpb1lTLket6kG1YNk4eDn/MKALKlTmoZC7mYy5O0VZ7gb+RwK88uZSHql4x9tjAw
N+NFasTSRzL/mRzZ9zQmGw1xb+L5I+ADvQazSAkA87rEntc16DP3qXoElJoJN5Qz
nyGtUHyWRP6Masraz/PMNb95DX/CfQKNdG5aqEBr3J5veZ5NNNhtG8K0y4CfG1CA
VfXapm2cBR6oJdMmxFpJD6tnARYJBewWLqpHxHaEt/EWnDMIr40gA4A2sHd3WKFk
tq/NJK7BsXcuzhpOOC7fa6om/8Oxt/ovjvavBMZRIUgzcDOkS/BbyJ4K9QLE7DoS
J7YP10l2Ay7qHaGrTzhb9ObH8uCEpDt8I1W4E1ZO6q3WsqDAfcZo48F2MyC3Gqfi
KrscQUQLe1ALsybrZdGZDrbmsRWpJQLEFqyo/A9qzKkLBWnOpVRkuYjmBvKVwNjP
0x60JvD1jcGicz/qfTrkIkTMqGVkUyGMNJ8bF/VlZPSQCz2sLGZJEpzMAQJswz1s
HVucr82DMeKZZBnfnyfHGFkXfds3YaxIK0YuHjvFMb+j3CQ5hC8qM1OYgaOSuz3Q
3QZpAyZsE1iKLCubDycFqeyKsseKrppIYl9ToPzDdZHGuwQWjtbUHWULJeescKdE
SNKNIGyMhCOJXKFmQKHhGIun3mCBjy1OZfzH+nCqQonLWdGm6CRL+HdiyNhgC8mf
rNqhM4Ig0h1DpG0gICPgfSdmA71q2TVgAz0vAZEWGLyvOh6ou9WYtS2dfav0VmgS
G4dRqhGtsRYguJHR1KuCLWKiDqC8MAVp1qR0oXIxXWYt5RuayjnbSaVLWEFPOPTg
uxf/D82/77kkQVcPifztLHX9Or7ZB5LN3xNi8ycSHfW/tCBVB/GcHqQXSxDJCQHP
VOqZkUrPBamqmuraI2ngcQ==
`pragma protect end_protected
