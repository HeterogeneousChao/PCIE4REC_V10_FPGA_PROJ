// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:21 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MJ9vh4E+7laxXWD+KsX3Iexpu21hLy3tW6PwtMaIS/QW1PxS4lb41yZmvYj0VjZp
dM3rgIHq1QvxjUJycxheqCL7AF5TkpTQQEeNzzoFpQg5dlGRlM0uze43ZGjBT4Ca
rAZFPJ9sLL6kVpTT4MN3bRcw9DsA7ZZfojoNlaL5WEY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25664)
+rKKjRJVM1w4Ok5OpVTimcUI4V8cErgw4FwchcBKNHfLplWxiEoZGA0EFxkJnrrl
UyK9tQg+iimTTYBdBMX0ryUlEt9mWITnDWu5q9Ui5v+GYVlZNpW/b+jPez+aOaoj
rQ68eIZngwDy9ADZKfn3NzpVgF9twzZl0TbMylqU/r9GzrUOnBLXA5A2feNlFhv6
dEiV2EamVF2zREjrYJYO0nl8SPyJPSyQFl+XznfRwizy5QDVeuxaq9iACyko8B+7
HqmxxNV59ltfJqmFunpcgGNIlQ64R2YOcLcmCywJyYf5ZKOGXIpahrckXadqp3wx
OeF3DJcqkJlxa3CNJk52GZV5zrKsHAydf7WfR4uj4rQ1cKFyN7qf2jXyYnr6C3Jx
ygoJa1+P2Zw3pdvPPxnQcSdonZypK0nIVyRuWyw3hkQIEoXOuZlhw88dit2CTxQi
pFdC0m29X4Lwk4f4MHFq7HJWkIwv5fU7Eph1DuPG3Vdi5yb/wlupLqr9MfwBFXhH
rvkhWPVHeAy/Keu2I+IC7ojtUYacdvgFs8GwIhTG3wPxCE3BxsfeMQqQdg5raSRs
bmKosUScVSGVCmMgCITKNBl8f/uEJvGm7xCy0cTlnfuwi+xIz0PlIrl6CCYPFxfH
gejkrxVuYoM+9+3jA/xaUvwMT+f25mzzsN0NpqwycZMFLa13hfQ0IdCAuTyZ566G
806+7Gjs3E2fPF+KtFIX5uwROAHkbKgekFsRMPBiGPdOYZg5BmKTsLBrbaGMGxNK
cYq07lDvhIckT5nX+aeiwCTkVo7MEntPXZ8HZszlOYOwva0RfeJ3rc+lgUQW0z4N
pZ1ygpvbHXiGmBj7BV051N90KPP8hliRlmJcqvkkCiFGEMGLbdpxOb+++r3PWiw6
9lxTRPYg3MwzfPoM8JonOqhOkGmL6F75qjmGdl4hxKjiw6WjESchUdTQnfRXEj7g
JOYK927vTltlGo2anF7mXzW5RhWHRpkEcGCuf8lgrBTYsPxq7OWd/cBZjehUCDck
ffDfdJKaoUjQHjzTT7RQpIYsWstaM/MWkB4GbOAu+7EPW4lUqFklqC+ykQlcsT0X
CAGVgIEcRfe0g5PE+m5v/9UDJ69QOOSgtM9ehm7FiBauM+AHCr5cDHLg3WYVork2
C6fxPin+VwXt3VFX0+pyKvuOGWg2QNU0qI9c+rtiUd8tqkCvzcS2UbZDJjOTWOkE
deXuW9M1n4TgidlUfC42vA186mvdsjtte9XMrFy89L94JG0Lh+7CvPfO8iwUtt1F
aTPi8aKck9xp8egwAnnoS8973TsRQ1pzkELo/CdjTr+f+L9zwqDdbf/Znq55uVsa
jO04C/l3O+gQGeWaNTiy+89CId163N7VbDK+mqGnburhSMK1LYE+yOFp4waEM1Xv
uzM2fFn+0GZp1WlKvxzR24ndh/geV4dzSlv7BQ9Z7VTNQzdOgFBfMxShbwdZ9+0V
1iBN2aMkDoS84lG5MuASRILUnSc9rKyXHaulviqqHnt+vbEhBB+ipFvwYGnPIVHb
ivqxJFAdDtpHJ9G+R8sjeA/el23T4uLj527XxNSFA+URTHpSWK7zEG4j9DnPdIj2
GXF83x/28oVsmqqaplAroETZ2tZLglfvrGRosX8re5zO5oD5Uwe7BIZ1wmB6WSH/
0rm28d5Va3Fu1xKiyqy+AwGt838aRXXA4Vfs8ghOAGutSvymAdIcLyv8TaK4xH5b
nR0THjEGW5NaNCK9ujl0hAeLJGmVXmInse1/J+xiSziEkYMvcqji4miH7Q5/aGNs
ClXCFuOBvYfPCP2ufAYVOOH0LlWvlFYJIrSpDSgIx0cFWOW+8PLLHjdtX6BFOgeq
mW/2uSH5Rs4NSQjjWqgzKsNlOvfAx6tFWsM8DYN1084LO9S/O/9LRfLsBqQagHgU
iKADOVMCo96CX/aMYiuUJSUoO6qBY5e+6ok4oGoz90IMIDHjFT/MxCyLiQF+A6dM
Eybv/r7/w1NEjtNZN+dgFIPe+drqDiZOCpZHHr3/UXAIP0BAmpzd0bnxZBWpIVkO
qMF3ppBrVWaPdvjccih+yz2GEw+dkH9+8gka/meBXQm5M3Q2OE6u6LflsPdQ566z
iMS7d05eyKIEMYcamyno3PS3MJ82LNmEQn+omwQp47bVdO9nbymfqkIf8uxdBaKh
oMMOKdHUO5CL8CjEPAK+pMf1T9SAxw2RJ0GJf8w60k1KbM4M97eyEOwlqNmbzVq9
w/XrKI2o96J5bVtQit8dEADYxJi9eLemOJqhTFWgGT/YrpZqveOvUiHpEsPHTn0g
dK5YqhaMMmFJruP3Ssk2JbauPjErOUpwEfIeT5T+0g/4CbhmD6Ijz06Ekzmrv44H
8aomcapIcNfAI8ksVpB45cVAUWNwXywMZbdVUgwiDI9kHdVAifbJToDMGfb3BE+D
QyE4/kBpatxoiK8ckb1DhJkjuAmAKHKH2cicYC9IkT9k1Cpd4BjZVBMUlvZvU/Vo
TIGtzKpyFltE5j8e5wuww4TRycG0/VMvY3JqCnSNRo1jNP/ZZvcj2/cU1nVELits
XGkCX+TwcMyClbzAHJrOgTHvRkcPigqPx2ymm9tvfPmRs5CmteERVBds+7CJ2l9K
yig2JTg8C9as6TNUs+8eBYS4yfOClmHxpjJkUh1JwhgmDhOO63UCTqilH8kVs40K
7yhQmoyEklFRUmXr6mK/5dDmTw6nagUrfZGj/GEAq7mdWUITK8By8F4QPBW+Styu
81IAg/yGhc9AHed11IRZl5ikplAE460y0Ey3sE/FUpbi/d9wKlYwM10/k5qm65Re
8i3nekzX8dTiUBKVxiqxFTfGdU4hvm5qLsn1zbbXBGQQsiVR+Otet/rSuAKzfLkM
D8h1ykPkN5EFT7jXYNniKxEnjnjAk9spliFRZXvCcvy0mEMOwsKZQrBdS1w/mLgR
D2mVHa6JkbRHkKK/dQuZUoFGrAhAv5HnMOS+GggdhVE2tin+fsHxf3pd/Uui6DPe
1X3AuetsbKpajHxFZ/cyoS+WAtrGVDYAdYjZG73gYB9h8oFwIj0W8OgQSK7Il6yp
3qComF1dVrpUy/KGCAAVxOYJAMCXdFRMgZM4Bd5D8q9EmbUVavsheEW7UWG+FGUN
KsNeSVkdn4+s6TsDatg+TVhzzF+GDWWr8QTagWCsteh7723uaR+fxsU0J1ycWnfR
4inv6T9c9/UISIAVrRnjVrllnlMk3SeEWOr7c5NxFxWS1NBDghDPK+r1WofWYW9k
ntU+87rV808oIkWpbD7vpj8fULHWIcP54Nc4sCKIzVmI5WKLfZcIrz0EcbVxrWt5
8vrFkIetwBY3VOItKOxMEzC9ViYG4JOicuy/sJxrruAB4ssR87lO0YHeKoIDG9ot
uPGc7dx6JYSW9sy8k1jpbYl/dF8tbg+KnDXYOE9ixkpAVRmV9SJXW0iakgu/6ay/
f5Rq6IZNj2OC2+TfS/KBAuSZNr4bE+R64p/LhVBezhL6BuoDBgLMLFM3njwHxy8d
4/J/bW0lexu9JA+TauekUt3LuO9XX4WOJPJpE/hAaSo2qO8ClP1bIosOiFoWu5Cv
2lgviBvQcc4/hvolaIkcuMOmfRkoPQ2NTlHOHR3HCb7eZbtbcZXIvZjc0x2OuvPv
OqqdJzZX55sqbRteZSnFZjDfzyXOo5EoiNiGiMCAZyBd8GQP0c6cLHzsNZUrAMLK
eAfL84E2gcP87L6NXqihGKQbO6j4+Q8CaqDhePiNulFtimJuRzLp3x6NS+zIIPmi
AIuGiNZWr89N7uNPFWt0QnYav1VGrbMltJHxZfjZp9LqAc+aKhuX3OpxBx0hesn6
C9fBQtPPu0Zjovl/q/QKnB5zbyDsWvyHsX4M+L3WGogNXoxIMDl0lts22HZFDORS
rOdqjwcppn2D8pICSpfjiHGaACuxjFUiJSkM1j8Dj34IYuECTReCG+iC6AmnPmuF
8LfSGMGQGFG/QhzS1ue0nI7lAExO9rOmr6fcF6D0lPRPWSXIuroSVvOE9WOoj9F4
YPIqFPA9mm8APFrVdkr4Xi49KmI1xBTVIuIJzloUmtrl9COL/Mpjs5o4u8lLPh6h
wl8cLTlvSGLu4Oo2V8l0FS99z8tvKIK7MTOXwbsME3DSOq9aUVWB22yi3WCbAsFD
Qf1rurHcJ6w6h0yADsH2GgUM6+IJ5WBzwlVXylsIi56oCe81ua0zJVMpmPDLdD0w
FdVP+mf94yvocGO6fDu53iFa+Q6VetUu5QQwgz7QvbcNXlh+3l9MYOBmuRhQ3fIK
pKd1InVk+mnwX/7xufOcUh2pnVuNu43FO7ezbblSYh86l1GxSME/i4M7zR2ISYnC
MhpRi4iZuMd5hrwh9wx2qEje74LdhDF0GdNtgaJhwkmS3dwCbE9VJF2XcFFLHQPA
DqWhHa0D7X5qKuoKYlFQF7A9uNryPUkjDBUt1BaNNvubtlspQECXnStWvTTyVlQ2
K81J118x/529/TNpvP9GX83AOHoR8LqXGdFfBTUXrhfVQ3Pq5S2t3Cl6nHQU0bUS
0gEm6dDoqzbrwda8ergNRVkj8UJ4DuyTjSYtie+P/U+zIxBkRvWk6JBaKnETTDJV
ts4PIEqdlWTrD/n+ryVUv6Sqs29btyeWDTrXqkUEDSPRxhWSU68BrHcTjO/FmsBH
ud3Epd2I4OcqCbKIsQBNmLXsiHBJp3wTPbP44lQkIdFWMV5EPPENHGJ6pCy4j0QU
E/CdgrAJVexe0JKLMHVbjBlS3Byn/cTG0AkTQtYPd7Jf9DK6cq0M+hN6Zq/UMm1d
Pe13jyyJn3an+sSYySqVl3C6DmE8fqe+kkaDxZx4SZjuIL8vmzC653LG1j+3MF/Z
LzAdfIsf8z+cH9W8WD29XuTUzQlBITFHPfLGBIeg7pUPWcBXexQtNdLp3Kx56iq9
9QUgDfTnUTlPkfbkdZkIvDgCp7M51qhnF7SMlKKhyClbeHDxsBZuZT1ewdD3PJkv
jWn1boOIQNKSVTYcM/BKN3qFKIklnrGcK349ap5j3ySUzOkY8DGO+/jgodita9kl
vGuxiuhxW98UgDRBNuH8raFOgyNlbmSdq0vyQuT/BU1GXsGN8f7swtW9osLPaJQ5
ijYcMetbQ2gS3fw/TMToAVrUeviDBaQDDBChtYk8SFTWO5LQupvZSK4e9G85ZpeK
P2Be31yNBVK8cAw/qEpqX9xJApRCXnS1Tugjjs+DttJJAK5T1dr33XZY6POQJ4De
iaWoavR/Qb3pbIZP8zuvwWkHvvevjAoMwkkStGzFXkWbUyly6qQePx4dsJnpV5Rz
BvzyyNSIAIK4diZPqciUMOVGDF84lO25nSLtu01OJgfxoAZbVHqqu50LTWHYQuc5
Pq9ehPfsqWtW4TjBvYEKrObhyVfoJQ2ckrzawAmmuYEo0SliT0g2rVj8iEXMFU8r
QE7GXOJgHNTWCU1m6G2qoM6WoMrpsqO8Nz1T92qTr1a+lnADaz3ASgPxUukN/9BT
NGIRsj/AGLiclQ+Th0jiaB3AwryMuM59CgLZgB5l+Z7bDitseroxEdZLyB9wE1N4
u9PB6xjl1fNHWtczZ257LdWYPMAFI20n+xgcmqTHGNoXxOi6fCv+9WDxPtfBenZ1
UU4CkFRX5FJD3/6rn/BFGG5D7CjPxZo/P6pTnIcGIS4TxOUEggr9WgvDQtOZ22sV
LqSN5SvpmFjSPhTXArnI+nR4eo6Sk7yAef1Xh6CtukKWJBqaEbBYGOQZFb9xsSNo
4DvUQ696fmbRDQDcZZ/I3QMLT2w8y8GpSiVPcjhuGCFiRt9Q9IQeqkwPwyhhSNcS
bx9+K4M5Nh1rk0E/zHX8L523iJf0WczzFr3P36g3pDf4CgFdA4LEOT8GDvvbb+uZ
1Sv9yvUy06sFQARV2fqyvR1EfX4pml8M01PT8HjfC/NY1WiCKbqY6p6HTC/PTDus
AW0SnKHbn8dEtzasXyBufEyCgPLijs61EGJlrF0Qkg7Q7aP9J2xvtpTdPVYGrLUh
Lg6/bfb/jgjkRUguwUFqfg31UH2SsNhCfVPuLJ7jDBp+dByRnQXcw5pcKapzC+eu
gAejadzUnhK6E25J8u83gABKMVKySeAar4zj2waFnYQTwh/74KAcULCNcQk6M1Xz
SgY6qOLyJJVqQ6NXI/CEHAM9YkpDuE0M+7jj6nqbDkTW2LPDZSxkNoQPMR2hVqex
eNMCJX9fwm0unuuHPKDO7G3MtLHEw0gsLln04k9+NNaufGet4fVvEuG0Dc9HO51T
79cIlhDWUjn73W/tY4mBjQ+LVREQIX1HJKImpPZyY5vNFWnuidur3TH091Ra8ijp
WwuU28+xuBnvVbjib9uzMTc3i7OB0N2FEff+WeshYxO+APVMlQ+R2FLudACvVa3l
IdT4WkWgpHi0WC5ocEiwO/0lvoSO1Mng8O5aLtXGBD6OQ4KWMNt0FIBBTTL3r07F
0IpIorTU0QeKujxd9lowfXt4bmGZCCd79l0EXOY7GX7caiMdz9O9XX5J7poGDPuL
T6Eb0/M1jdzp8q2DtmMPbg4HtkaqAa7zaYonnF972DJLZ1FmjHE+BwxJq7EuTNBu
2sSZuCFzhCrfCq8+zcW1KhVWry1K+ocd96X/2o6UAn2ULyDZSVQHNWHdFiRGicXv
yIyUwzUbmILLZjGGNs3MH9bBHcZqT8CppscpaW844zTwABjMBFnOoPSoZHxgvoyy
0bCuVW97PepRHa/JJgiKLBlQjTcjvAt/rABBBQpab9W9QtIaP91Z2KhIMIXctp8s
kmA6mDLxuApmcS9pE4kiptjNFgiuvuGTw2Y//obUhkdRE7q6rBBuw5pzxhNaB5u3
HG7Hs2KbyK9CxjrS7lwtjxXPmZAZWljLbzQxXeVio8HyFIh3W/CN9FebbxBcCg+G
xsIqDAN/Dyx5dqvrZfsmRi1dFHOIs6lMHVJOCrx8paEwEAKJA05MFd5BYVxVwjcs
W7C47qm7cxUL7Rxl3Ck1NpI+Dw6i+HejjP1TlAqyNL4F7rmibfuc6ihUNH/wdJN+
W/63/rSa25xvokPI+GoQx2SpToVK1hw6+8HdIUosCyu87Gcf9opL9L6W7kXhSIdD
9fCC76kj5CpadDVqJ4PxxM4P6u2cYh5xpnYFNZ62U1zQZJ53Z7NpbuLXVy01nuOX
nG9xYtQeeiYWM/x92mELjSTEx4GMYJd8HqP+3gNh6rAcqeTGW1ZHlt5gjVRUiqZx
4isIadlr+CfILFSIN7UH9Rq9lSUpaSf9WAAK1yr+59qHY/VcQrK6NTA7si/FRL6M
Wf7xGh4YIFc3WlgFXefBHeLbR09VEpEyzQP3C7mb97scj7Kgirs2BXh9iHzWwuHj
XB6KuG/B0lT6I3PM7kuNAVrkI9LjA43P+/L8CY1Ji6t3QkyMLlDu4K3QCLB3OtDw
e3V5hE3qJWUTYnCdpBKK1/dMB9h7UvKOnqndvYAenNA4loXBEKqaHQtyDIv7ko/2
fXnzaQVcEaNSGE/6MpFDLC0BiPUMLHdE8snrNMaqUQIh+0sKO9m5C26lXOKTPt3q
qChNrieTaDaTY5WKIV/MRYpLyczHeiV4QSKNwZNLHgFYxfV3h+DFQQHNGhyVLW1U
/ges3akqp9uLxZytTBV/abWsyVh51vxS7uU7AjZqU/Zl7PCuZrUINEVqTqJgrzIP
l+O3dSleeSj9VvLyI589ggruIGAsCrMb39TMCgVETXuy3mBjFFz7fBwR3R4apNUr
lQimVnWOdFrHokqN0UaN7aaSbdXx8490dRNae99P28vrVNSsuLjY04Q5I4ZoF2y/
hOLu3HkRJNm0OhyIEJLTLEoae+hKfLnvGww7bpQJbGXH3o3TTIaryBLGpbDKXXQ1
+Su9/M5Ww/GqVJyKFRP6Qw6wNNc8PBT91sq9ztE2BKKEIzlSSZU0OpSf44QSqm0X
dVdAwNTppXMZ9rU/GsUe4Pt066fB3O1CmHkP2ewX5u9u61O2ZyeEu5hhehKrCMns
u1EzzygdZu6Or4DBu6a/BP4EoOUh1ADp8T1L76fTaZNCpld4PBVHf583MMLELGFS
YGx+GUr/LQoSJu1y9D1Y56Ga2D5MyY8J0WO7BNiYfC+niXI/tsQIUtfLrDrroDSK
fCbWcWn4v8NPHIHROBJ3kDD+bbdB9X7M9q7c7B/OX1mkUvPIxgazmH/E2FilNPLU
WZyORc5Glx6PwSs5WvUSZkNHdkNhpKsAKC9neDm7rFPV39FSP38A85r3CH5mJq0z
NCO1WDqHHkW5DZykKG3iVCr2lUdqVQ9AoQaSYiVpo34sVO8WkqneVxuKLoapR5w2
afyP2ju4Qa055WeRE1CHF4oxMCyR4r2F5Ss5eRdUpgIhqo9WwDSWnXIIz/b8GgZs
3uq5Cm5GJGSG1ElvibzSmFAK/whUFuBNeW2ezx9HLxKT0geLtcXmrLZUebmZTKe9
5pA+yOeSvWpJdqkvpP6J+9lieiBCU9iJLg9JuTOyDORMhuAwrxKO3kmRKNDXHEbs
Kmmt3OQTjMsN2ESSM/K/0uAviu+jRRDY80rH/0Ci0NvqyvajAnOhG4t+IwbZKS5R
OuRNkgSOYcXrYKtoMNbEHTlVfjSKLfE2ZHVwKWZcDyN3sRskvL1LLmuKD51jKHQU
rb6al2oIEFMNEYQd36BQkNOAXLfYdZAY8x611D9we9jBemrx1os1tbEEeA+L5Ji7
dfJovKnnJAL8vUPGJlJ6kRpTk3EsT7n9mi8RF1dA6230Fez9Or+U3REpLjgbhoXJ
WiOyThS8cMwCmqWKoysMfh1sLCBNOT5bY3hTrIp+HPqOGy69gMG6Htue4wWtSd3G
U4Yk9fVBWal7TEmxgosCDeTPHvRZW2tnZuZUEpePVOQFYSlenL+zrx+fBFaGrN5P
ysvZx3HtiC5HfSPcg/v3j7bu+kW7h/nzH3XKKPQNPB5qqbhlouAInBRU5NC8XIGV
LAnJFx+r7p2tiY+cdeQp/Ut9NWz5fl6enzqQxKIm0/0LEHwhWrSngdBw7OKa3mlw
45ecy0jLvR927iLhSz7MMIkU4EQBr/kfGQa4ndTIUB/VR84xC63v5I/DMb4dUQqG
OqjmH/1HwsIXZUfjVX4iAoEUnjvo2zOLhHzA6nRSmopnWPPP0qBct3TCkKvczDLw
XWayXfELiTIjd19KeJ2l5K4WfoxLpac8eB3d45bkpmA9odvnVk/6O4Ekr49+Skr/
2laQdWZKSwOttsgZzD5JUc+eiDYnlq5K1NVP+C0v7ue33aKSG8x0iK8oC93CRd7T
18N6JH4Gr1uaF3VA1qbIza0CsYpQAgDIOthfoFlLA8vQ3//1dTz6buGm14qDVnbL
OXWnj3wVpAjbG9R97GTjbnG5wo0b5Qa0D2FsK4uqv7Fbd3yKo2FR8WBoEnzfTALT
Zm1switzahksvC/0iHlZJwM+xK2+7mUcNHllgc3oX/QfeVmU9d60JYkEfstMDmw1
i8YOHjDOvOqI7hCDm8rFJ/mGzcFGOdoaUe6jTvCI7yXfyXMqrdMUG0f7/vf4RhbG
14HojVgS17xz/5wqowVtBlOr+8yQKJDNNT1j9B+7zGQpESwZUCuQIC/YT30YP+/N
lg0mVqAG1xYdUZrZ3CcUHQoN4D4Fb15nzrDZ8lmj+DTEzCXVlFIniJb1mrXpMFBW
OtWvetnaq1Sh3TfhDCDZ5Wo5yBevTVVflP6NjAVrCpzNcaVGm4G/KB/cLQ/1KVar
qAvVSxqJuOooBjkhMrpF4sGvcNaI0xqrLCNcX7pcuKdtgimDD3k7/KvJ1HQ/u9CY
Rj2z9W1DXQWPKSE2TVmB9w+LDqzeYgH2OLLBdyICLlagikOVBwTjOlUv1PFEFzVd
r17KAkTBK0hEVtdyKRZ5YcPoeouBq1nG0SqVK81GnVdF0CRqifscKvuKz/zIy07g
JKNXkU+ewf+nyEKaopNpGeVaoN0JGCAhdFQkNzWvV38fRz8X2drnO+Nc5ZBckF8B
42J8SZ0SUMpFYt76AlhWdrKFpokXuS9UALC0Js6BnOVZqayvVvqKkfvuDPmg926o
L38JERzWfXyZ4e3HKpx2RQ7zL0M715SJYQzCkCFgHkV0a1vPqvRuT4odL4DR4u1j
9NBCwI2AkowhP5Z5snhBZEHdZuQewcjXZhIGzCNz9Cma7HocVvuj4K7xA565EAnA
d1Or7/hD3fCDrZv40pX9iVtf3LwyEtYbX303IwIJgHK+YYu81B15ESJ1Zg0bTP1O
E1YbveeR0ebsBy23nFNs58Owbi9fWyhLpPcEYnJoBQKCTcwiyPrVA/vk03q/lfh9
GR3kSppyPy/0It7ngHxh+58cbmoCI0lDeXrrTVson6irLnnY4WctFXv9cvUbFOG1
6GLnykLJzo4v6UG+roamBceyOXCQiEn+jQHY2Ja7IyZQUICQQoSPevVJapVGQutn
spskuFomsP/OXoDCKA8UMG68UMxNwXgHOMzW05xj4AXRcIH00G5HN/saMa1o44DU
XBlZo6btYi3nlHeBLYyGiXdCzQQEkdA+eK2OcNzC0PqXlQ3+yxJgHH5rdtRKu2uO
60YZyzg8wN0FKUBALye/QXX7DIjNJwuLxda+AZkR1HazXvbh1TCKWv9SHmucf6BZ
I4DZyITqUholqFjh4BlzMn590z9Ye/6oGAzkTtM+YyEgeY0dnTu8d3o20LNPDMwC
FU2IG9NNamRr1YVPd8yMrqvdbrsHF0aQiIFb5OpYrDoVq+5tBJY17RBgoXfzQujP
txv6TLk8X1J5KvididhNlwIkNdKYCNbLdgr2I9MPJU2yBbDLx4hpkBlNT3GIFdaB
8vwU5Lewc9iE/sbwLWn4t2Po/7tns5tj03wDtCRd4SoSAhfIQt1rkecRBLfF6v+6
W0STSqNzjqRKl6dxwwYYUvSq9LAHheA1UK49naYlV5Egui/E/bMy9Wmee1tMTaiB
3i1TTO9OMwA6DjShqE1kDOta9IwGGisku1IG/riV8aqhsp4bHTejP8PmBDjObj4n
7pj0ADKzD+WA2pO6O5mzcyWHdpLd6sfd9YFhIwIJvpRKFDMgmtZsNVq3F2q6lQHW
o6UbBHEvIJRRGQrhFn0aWsaWdSKnLqVM0HjI1hfNUINJvbll0G8QfuEnuFcfGbjW
y5hQPG9djRFkfcd5SrzOLkb+D3a5l/eRJ6SXWGkvRYs/h0tFth0r8eqrrvvcvEgm
uXdT9IxbxVbpthkgJa/1fW+4BQeOYS8ISRs5wlkoizC0hJikGUhxEdnmyc2VzVVt
pzlEdi9zXIZ/4aezhSLwAhZuGxNZTc1+e3Gnht437pyzp76rfJ53jB19bHFGGhpZ
qJS5dMo0JG705BTOaOHO1Rs7agGnDgejqMT0muYWaSCvkrclqiPDS4Ds198fThGt
BmSrKP98w/A1IOERDGFj+dAxdlSGqjs2o4UmvEwU0pczE2CO3GMhe5hcrfKFasBJ
RpTqvzzmBjfDKHhtBBR8cWPUMk5RU4ION2pqsfzaL8qAsZWDCM6ZbxmqSNgWRlOo
QCGUS0YVJbzoFkoiAp+k7AsK+tcE/I1edfw7iz92Os+9bLSVuBFt4Qia/hlW+m3P
UUdvHjn0QPWiMYLmXZiJvS+NJ78bZRFHk93u9KTXQhqDJdv3EnwlYvJTZWn8cNuu
8PSDJaGSEvGGLxwlQCrB3pX+nAwsoSldEv9rmkctJN9cUyl04v+2489qE+dNISRF
B1PWvDx+lAgADpol6mX3MEv31L+2h6otdaQJ5NknKwnLd1hqpz0x/dheoJhsvN5C
bZgnECaOwzDE0bm8km9xSsCcZkEKX9FOygtVbr9/MLOX5j/eb+/QYi7joWGXweDF
j6ACuuyS2WDeRbQPUHvIgHR9VQSrD0qwvpnX+SLBOkzdjKqxzED58Iy1p28ixB6p
aBKe8urwLOlFvaffiHT7OLOE/f/4EYninqE1GruGkai6ysqDszxnbf5n5hx81jrj
kGDIZs5qn4o+Kz+1Dv3ngnsM77fEOE9Un9IX+zoMhpc0vPCht5iplKRI1SNm7Uj2
/q84IM55luYtH+ov0Ek9jBVfQrjhh/njWjq3Q05S8TF3+tk3RdrRcOZ9575zpX91
t03shhlsCh9MzdhJOwKHwekRvk9kyx+HHgFBU8h+RjbFtrN8MwppXxusZHUlEtgg
an83CNEDxY966c/ir/r7ETO6fnHLBcHOYdjt9u5fr8g74QCORpvDk/Wo1DgWng1v
yPF1vHZMwFLUB7L00JvbZ7HAM+lhFzKIBslyHqpcf6zIgsZGLKQGdKn9sakDGSIl
jxcY6Zs1tisKcNMK/QkX78t9FamKQF7KqNEwpX9DktAaTS6HS6JDGsXpai/BNKkw
xHwmD5pw5ZYhlNmz6adHnHuMg60cs5kDAN0oiGkZ5vVdeOZ+mOvK+vIrwNgsLTH1
z87PcMtm+i6tgGcuWHjgLRvHnOQmLlHZpcrB+Rm5A1jbz1RyJt/1lAU5cqbhli2v
gvRVWHNdS1OFPyhePMLkD2ottciLjLAxFq1DKSChnypIlyOoaoEjBX+tg6RD1Lyw
83Q2HwzbkQgrG4jXBBcJQGtR/zDOHUkoi5ElFNIZEwWrHeCrkJdzAznb/8MT3W9b
pFK6uwW3ahBKG1GtfjqgEb0o/KWM9GDtj9xECh14qv67rIRdG6HkbWsV2N5NEYE7
F7Tr3SidGNq/BLAwn08ulGooRojQrj3IC+BIY0AAyBiJZq9y68WXneOqVAjbQJmq
9HU7wN70U+6IlL2zIM4uByuIiYMJwrLoQTf4IqFXFCivUgis5uaKzEL6YyhuS/tF
CW9PNisadgymhWyPMFbygAVMw9FFYz8zl/yni5evJeuMgW5goVQ6ErG+hyjQZr3L
gxDKcTPmO8fRKPaU53cdbrtK1wKFGSbiYlj29gwd2mB9qPGrNYHjuoXGjbXybW7Z
UiNsVGLvl/vCulSqODmQvhil0yRnCQzS4SkUz0Vfw7xt8atT7eoMBwZKls5FgQ+R
4C2KG0yYxj17js7NLAumSSf2M4+Rbsq/cOSATjkr6B3ZaLwuAZSqeejofpojKlHn
1xTBCwuUb/Xt99Vv+4x7tk0rLKF3Jcja6vxQJyCAmZ0RB5IiPD3E1XYpvF0XJeHO
Fgi1rE7KvqXWQn8PcPEtPlo4/MokBtLjdu9SqmaYBIMoAeoR+kU5Qr+wNhOIfZvY
TimFkr73Uvlh5L2Hi2BIE1+pb+Pbk+wWf5AwvoXnnJG3SbtqTpoY93ucRhsRddQ9
5o+b53dVyYeRO+jnYQmeWqHWJOzzsoGkUwJ9NeNautYXTomGeVDNQVlQ3HJz5CoY
KJ6Ng+9qKlJ9XD1aoatyegh6o+fYcMeQgKFP2HSaBmdk3FZI155JULUhjgr6oU0F
G/9Wy4k+K3H+lA0NDa/OXHNoe2W4l42scZqcgUQq7jNE4i9ofLI1meJLi1ZTgeBe
pQeXqEmtGBTrbx9/Ryf3zKlqy24Ki0sf/zLGjDAys7LAgTiWu98zkhEhjcVTLuUc
bwOLJJR9b5B2uWnKWCsyhija9Oc28eHszQHp9wOY9LG6NxS/+H+D6se8qF0KN/Od
LhltaLQ8Fzy17j95ggpiBkR5mcdSCD5x/NsRQt51AmykmQfDre5kJ7zYylqhmmUk
922FTd45h4N/YUfVtWkBrdaMIQG8ZOd+3rqIqRdL1LaHHYRsI5iU/fGry+fQX36X
ug7hfdbmLQXB14aTm3JsUfXv8rzOCc64OYHdnyWVBdedsBvqP6jeoat+LfqTxrIP
cUKjJswpvEEr48YqJH33UTSWS9+glVG7ypR9nBqunf0baLMFsWJp+EtOSwwm6Zhz
/mK+6tEQyuArc3rup10uH+8Yp2wCmKT8Z2cKSzoCRwy2gAPIpuf9D6mdzRr3uUA8
5TNTW5WdR69tJSbkYvWZ1JATMVydXH4B1x7ae3rjZnTa04O62xbW6/JesdUmynQc
Mwxlw3hBEmZI2Vl1E3rQsO8KoiJe1tiFVogpUedibmszNhoa4pigXa5bl19TXlqY
W6n1bJchUtpKIkU3y7zmXEm8sYRwo7ujRmx9QYsB+zh++xjdBHLS6LuwNEejGrjj
1cwyrcKK4RPhaHv/8kJbAz2lYGaXbpGNTUgYLpfoLvfZ7xFptOJqT62Ny7IURhtt
HPg+SC9HB5ZHVeuLxjX2KmCogIyoOkLbF4+DX5muWlbY4g/6asfG/U7lht5L9MJV
mAxxkc2TLsjlgO0Om5qIhz4teWTTb8KBWvMbetUCXSN79OPww+CLScYqq4XcVhxX
TrGgJRXOsT8+Dp8Mx7DVJoLLdfyG3SCuW7bF2hS3ePMBLkXM6gUOFVnkOyx9+bKp
pcG4MzhvZzuOj4I5mnh9zNUH0JlHFZuNzvMxL9N+cDTTWlSeRGynpTQlszATnfBf
lH8c43x3Xzao6PME6BujbEgEvJZ6q5MDnlj5q+wY2reeDwrajPYyPbRmld2oSXzU
6cbkBAU5rG2iNTQAboA6VZNvps5X9RsDmLcrGNbuCkRhOyricbafHNT17145Ch7e
a87b/lzEobi9BO0Wsvo5IP/FN5CiXcwPGKhei0SrXHBOe3VOVCa9S+4KqpkKynCv
bT/ae0mfhQrCGq/Bf4TFpf12Bka0X8DQaBgA29D4QEVFfz4IngW4r59heM9bt0ba
YmnnWR0JsO4aHBmu/soO3tqDr9r2sw5N4ZCvYD3HkwpjnlVXVZKpEiHh7O8OABQy
lvHG9cZ3Tie5tMO5iH1KcbM+nY04mPDaUDtF6dalU19Kv3fouC1seFVHqx7F/h5l
D6xrjvA2/iJSnm/bJqC63JVHGd7G7vzew1Pa/kazqa5xi+suxbzg6BAV3LmxBPaM
gRP3TwkdQnnTEQ0ul2UKusQnLk40G/xNAbNxiP8wLoJrsXkkv/aFsIyo6BZwwUzb
NESCAg+Fh6wQgsNvN6De5ZfESQRPA0/D5x/zekROthStufQdme+6A5XijqvwQ+RM
REe3VHEO7P6Y0KWmXHW+6oSieMbMwg7JcG06quiOMOLZZWHmp+iLhjhwA/FWXoUj
nsvWN9RRq7edGsLO5Cg3HvR6qx1mzGy2nCyLF77Y0q9xVpoNzUtjO4fp2KJAsJsJ
gXzlnckTjeu7d3xFYvVSBC0gmse7jVZiVsxA/dRDCSLsUvgqOestffavfHGpB/kQ
Ai9/lQpcKGBEU3UNqFVI6WMLnApKSVw+vSevsqK3HPKIvE4QeRJrCBE6xIsk591I
HdjAruDbwYKBxll/6Cg/QN6Zco4Lo/Rx8eU/PdS8Ga53DjYXbToOyV/2spR8pNZ0
hAGoFtTIvWH2nwXuuVJFrH94TzdkKa91C0t35PtsIrlG2wHqqWb/pZCahCVwMGrw
ag4oiWKkKclC08FCc9Xao+DyCxGo5TLZJZaNs8pQRjFOvEKC7/sDPyLmRLrc+oig
uHV7D6dRArv9sPLVcX8Us9GyeU1YVUKWegJ/oAJC+zY/VR4IyLIMl1sO3LtTe2O0
VSjbRi7yRoJDNg87f3z/mWYCoYqToABP04b5/waAGvbgdqHQDnFGZLLM2PD2h6/n
v4adqV7CWTN2oHNkNgcZ8UsLB7XSDy4fIQHzURKo+HdBbUgJCLHlvZ+kQD7FVuPQ
lMriLXSa6UxpD4FzI4sBNprW/QyuOi+miuoPS/j8518hnlZR7jiSrV1O/S1ojmyn
V/giQ27fjXDNTAfAJ29XnwKPfWhEbPsHN6c5W5EodCZ4PYcwro5ZxN7r6y9hfgkc
AYruTF0hwcBVfmxwkHKiyIUtd8drs7lvZAuK6pT9MCS8Z+zvYs9KRfnds2oVloHu
mcVCSrlOcGYaPzeHuzEaQgHDL4Vc4Hch9dChyc6+Yb0MqI/pUUOQC7AugPly6qg1
/J2fVukaa1bX04/7yPVLSY4H4CicIyAH4jC7Wk7uehbV24Hl3bUN8eEbQgxhX17G
zZ/S6HEdLbjewmUp9zCx7sD/JEWJrUtrg+zKI6mbbytuldzfTk8UgRpTV+HzKM+A
Gmzr9sn+g+P1qICDLCRFucjDioKWdzP3z9gRCi/sTQtADA2NouksadimxY8L7aJR
XCZhOBFHQHpvHy+eKY85YhwIIvuupnh1SUpBLZT1SSbmcZHAfveU6fxNdBe2cf35
dXwEAAS3mo13E0eZTc7kA4QhyRf6WZpitu5mZwyoUVlI99ZUFAOD/50muSUx8Y4q
9AfQQ8L7jvkzs/OxyXqxqFyVsTFSUrG4SAqGa+aXCUocYDTEATSXY48Gq6mb5R+s
MAm2+JvmvxjY/lYqoO9jCwsWYwTUdg7iWpzfKfTDUbIbW8wBaYbWeNfUOQ0bxPHC
TiHhHk4Woujc120X9J0B7dJsCco9kCtl6wCYhKMwX3E+cDvHmCQEFDAnXoSp/3cC
ZdQdWeLmE07gMS+AU5ovE/yE54tG8QYE0qs/pBbStHtB/mqEAZunCpFczEYZSOZj
IG83I2Ho94W/70aGD6B7b1+JWGzIjZUwrLsHVpOA4hOJc4pHiABPXZHLkEbsJNss
AZROyG5SbY5CwRtEDpvIZV3VSh/yes73rw/n+ggWo/Shj19LF6DEPElJFlUXiJTP
2Yhk4SYTQtDLEWGslRNGuTzKn1ew21nxJegC6uiQFRUxShKBVIhsLCyVWnkNuO7U
XqiA+7C1F9hrgsHNCRyzTv2RX53JPZsDUdprulhZPda3oRp/S9cy9kj92rbPeZ9a
AZSeRP5Gw6ns9pYypwKGGiPLdh0O3FPAMCtpDSP+56sa+cAW2JEebSTouM7/fF7x
t4Rhf0ucPkiAm0kNJeN/+MI5RIl2pRYwsUmS6SUts9XNK6lgBahLabP31PB37/vS
T0aD8lrMTbiww2CWk6rfsgTO8HRuLV0nBqxJctJvH7HihKTM0ENASwvPfjXFGHKA
3i7wOOzCMmaH+z8UKzbCY3lnDMQ3yDRzSxZ1ep9FFTDthNIje1ekO3t1VsqKJog4
GSS2xIgX7HJGjk3t4m9mpNRD8Ih4jEXUPzHTgGXFDNSzxMNet5PwRQjnbneaBpV5
WRYkYgMyeA5O11qj8oJaMKNg3vsQ07v9ArgfWCU6G/NSMGpqcF2jUTFluQ1NzA0R
fskKQxbSJjn6sJ8UKwLQEOX4uF3ZF0/1IYahnFBwVr8axwxdYRfK/qlKnhTd97NW
G0mxKBfQh0mjky911rRR3+nyK13Epc3AEhxWW/CN81qWXUQnjw2FG4fKQCIlh5y1
GBUDbMUvvC1E5fueXZTVkr/xrNesO+DBFo1V1SIa1hehI9t2P2PwGQRebcDQkGVm
2GkaeYPkFU8YBGtIfCwq6kWh8h/KLeRW+0vo9CgnlSP32B7onUvOvX5EYWCNQz0i
KNzw3BTYunRIqyzVI6E8SSH3kK01z1ohuGDtpNykWdqiue66JlacO5hi+/O+n75t
4VmMX3ZjYMakLayFklGLbRgsCXMi+MVgZol7L2wwWcs3ss4ScjibC7pDZaKjid8Z
cgmKIIcWiHUfmd7p2Mx6lgTvLz1wnGkFOJ2L2rkxfmV3dR1pFU4yiZSwU0XxDkbS
anCI9ozPfEx9mMCZjrVtEOs6wECO1OuN0HJaUg39h/Pk6AG2G8ij+XdZjqEbFZlB
x09Rg4sm9Cg46eFajB7YJLIuBYiQltyI5+EO8ERxK9OWYib1M1V3sArzi0wnY9Gb
faX0F2/dHrhEQb/lyfi+oO15cve8e9wVtNIucNUrXuYNarVMvAU7oJIo072/gc7N
nfdjBRp0tDf49tOXJM8dKc57Jmv60iC3g0dDDZOEfuh1+9ZsQNUuvcy27S/HU/VK
9bib5LPHG1HXpdqNVlEPuMvk1AnbWznaoREMg5jUEEy8B+c2nLKBne9lBQ41ZjtB
QcIUD1j+05xeXfgl+SpanBlQSaaBDN0qL+GYD1ExWLsubOkdC0s70YWDrPHVTSZJ
URfmR0QHSc6P2j6IYDfShAOItxFh2ZH3/jN8FcnESSGMBWA7akahxpSgCh/56pLT
9xsOF/dSq1q+oDmaskvm0M5id6dzlY4Ch6pUNKW2BxmMqBJ0kQnkxE2RIVaqGH2a
6jCW8sPkCIksK5IWTZt9VwWpEasdSGEk2my/A2BIiF0nsBlSvSaqJG4ueW6ZGqN/
jVSa8Wy3lIYo1fPJM6ZMGWekbpMULokznQD4DaPTGP2wDRAoSwq0lDGzoOn3Rkvv
GKot00qUr3UbY1YFJcAHXOW0qDb8LxW+XQ10rlYXZvnRN9u6OKE3ciqQkK1eIOwD
RvjmyeLz8VpOjRbRaau3c9mOHEhUMNo8Vx0TQgm9K6nVN1JwvaNR2hlhAtwssw5E
zolVa4joGFB3JR2LtmBpQIMsJXCNUtw9u3ALi7sypReaMXAOVAlaJmIqxBvWP1i+
f2D22u2hZhIEpzAXh7ghSH0jfPrSJuFpJ/+RJzh6n9OrYfcDnyUJWpx/Bn95b/d2
eec+tO+/nHTbFqXJY+EF9cO/0wfI4Z4Gf4WfYUt2yCOFhONuk/A2hhVOqS2x8Jdb
2jpLT1P+aH0ywlhtSrcui7E7YC//arKDqvEzy2Usmomb0eMwr4CzGkQXLf0y5v+y
yfC4ZStU/bfyVfwJD+TX8Bu2MM2aq/r+ed8xS+LWw51FmFz68xq5T5d12/z9H5pH
lOxt8LyUp+EYrymL6PeXSgZFAgtcWwectmE5Lms/f9kH/JU+p3hJd0wFoUfjBwug
kq8f+SF1WkWOQNHdbXEC/tL6IaR+HkGitodzVTHD7llP6ptwhl4+N0zRtXOP77qt
s5EHCvmUEfZUecOdh01zHzwuRy5gD2aq9A52ieOpqfEvBoA6yQo45jzNTx/80U+r
rb5krOmCuFSycVecyqg0rQlndGWS66PBAcHxLTsT9Kix54oS9I+gsy1ZiKk7+qfL
ZgWWL31stOq/Ayjr6PAtTET/rb2/1CSPenFrgC9gh1+6TtEOILpo13BeBLTXbDgm
X4ipMU/S1cxPMnLeLvrTh+qTJyIVudcAXKB7D1SOT2Dnk4gx3wr+A0B8M2gsWLyc
/iL+2TmhiJQ+6tco6s/lUIpbSMmt05H0JOIlD8dZ2q7rm+EP75WoyjstwQEP6uAX
LOPV1NPT2axIruV9pDo+imck39YexCsVmQALIMMRUOVB3msq6TcGB8vb42fgMMaG
CSiZGeiC9V3uuignOW5vgh65shdPzfpJYQBgfIpWRuRjkdpKM0Xn5jcvbSHdXQQC
qYLPl9oWbhc+1PfqjogNJhxrkgpYyPGFxyPguWJ5neYSBveTTThh7Qs7HfaD87lX
w3F9CN7i6tiBDXij6gOeyeoby85RQSN43ITOrtwQGkBUfY2E9W9BxX0Xczs2FzIr
y7aar7UD1EIvbDDc2Zy/3uEn495NuY55ayJPfPtAAEtLt1caGmZQtCIQBCzrzqeV
JHBm/384+6CMzOWsz/KFR+01+gcgeehIAY3ALrywrRdHclkU0pMn8HkVTAahe95Z
A1wo7vTi7qz66jMDEq77u0UJ+Oy8U9vVwefp0jvPtgHQZRRQ9U8Vgf+lslAhYn6C
vGLAFti4Auv8ZSqd/fDUFTEO0YxrH74FU4zphAOM0q0RDP+QOujNYOjMlYXJ1aGf
uu1rfNGA2F2xPksrPIIHVPbjaKsUDSsTBLXeyK6MRHdXENtXN2AvJTZKI4ch4SnA
b7EHdLlW4rzXMDFqCvj5Y4vgQf1Ro/795k+ppjNK9RNG8YEpMlhbnEZ66ci6pncd
kf2w3rGpVJ8s3ORR+3cLlp43ZJKFr/TceJGyIPmah89+sy+h22gD1T8zmzciWQhk
41mg+mb8XYVgQNC5fAL+FcCHQ6aJPYXPCNeemBs+Em1LEM1jGwdyq0j2n4nWEKT1
zs7gADZ4z8hwA5Y8ZdJOweyRBRdUU5zXYiFb2TW6AzJ9dE8l8EQz3KZH9ex0u51Y
PTjPx0bQs+nc5/NdOum6QfOz3QnSyCtR4Z443Hp73s8AxbdZXmyph8MgnBOCsCU9
XXES/qeCj+AdR3In/1g6asxLJ2oTwnLcCGlokgU3nGqVCRcL882NvcHxvfGzM5rd
SVcYFgUP6oPRT1l2r6VxMeh7IBACepINjnF6x64+ZVUkSbX+crGlCruUBXdvR7Df
jlrMlv2rQw7bkzvjfWRJGZqpn8+6bPZmbvorBB7tBluN3T1iy1vIgCDWzIM5qOgc
vyxwxy8yp3SjBvGvVdn75NZLVaV+Sq3FWtBtLshRU2OtVcWTIkqEh0tk5tBjwupu
E1HwLmAM/vOftcNJJTGOrNIuD6oDZp10K1TUm3e5IZ4xvzXmX5uz1abPxEYdRsnM
ZedRLNOJQJE9qS0i6v0TyAapyyASzQGiz/npGaD6MCvmysAz8vxJS1xnrZo3gA98
IOokxfVCPDcM2zcknTWmlfdizTOer31MMCNvb3VWPa00i11xitvZl68vUsyGSSys
vHNHG0w/waAMLATuxzhVfdWI/m8U/g2l0KxrL3i4bdLP8jQOk/a0msiYB5Olsbx9
BXPfPiV3Q1eZrj6ekjSm0o2kWovoBi7s9UU6am4ACAI0WiMF6pytYr4Oi2tmYbel
EXnwiRCGrT01lJZaF4aLQDzY7hL3Oq9+Dq+Q+Qt9Ew/ok3FJiiqOrllpKTRKHDRJ
9YnOCNZAIDb4Oga4FiMBJWavjt4si5m+QRqdEALkRltDW0jVJZ+K8vwV1/QLG+Dj
ML1vytyYAtpNp+xlYrjwDShOAj/oc1Q0pfC4cmXlfLugSTAVDKGFM3fKkuGg+iPL
jTzVjwfkERd4uwXGWm8GmzPRxWfkbfvqdO8dKW1PS1XEZ3DzzoFLGeoHdwJ3qGob
jWvlljRtHBGfZuzSug08fOqTPf6qpo7a6QIl/nXvqTarePrDmw8p9I3A6O4oZqZG
BJ3mlxFNpLP6SxvkmU+yUT6/fdjeILVtg1h+jUHuyBVLRLKSB53239fN3dWpJejr
b0M0T69ZssMmHByO/QU/A1Db5pjSCIO1MTBhdkBy1ztsO6ztzVwKNpe+fvPAg7SQ
jrOvJWnJTTt54wtAfTg3SNe/afIUr3J4WqEQaKbnx2EmdukiJMwanejkreAqw2pg
5t944suGSdil4bs2MPLE4GNQUuF3RnuvSsqArFBZuOh1GdPLLgYwrivr2K8huPWU
LrsC8q+Hr0SIVnQZuSeKfEJEilYSFlbzDl9ph4uq4+WLkXDskcd8XfgIHPYUnGGM
QkB7P8dF2tAYyA8TfhAi0dYxdpF3AuwMH838/kCUOuRfya0TYF8A4oNFzLcPMULu
QJ9sPjfHn4zLZFgwe8uL2RVhgQS2FU1+wkEod7XoyTTUilxDKUemPHq2LUqtU5iE
b+Gpe1UA9GfEoEkca26ScC4D77QjDQsHkZXxYpEuUpuDZAx53vNXp43TyyMigyiI
7i060DHuBwPWZlS7Klx1Mz/kr3IraNOsEQXLrcKb02o6OiftxZsjc+NpCXu2wIpF
d42snO34x6MYKsRjVQAsx/fRNXfxaWp3H651x9ywm2y04e/zcqd/PaxujT79oNiM
1GTB+vrpT0Sun9hT8nNEBARuwpJ7NUSBrWkcgW0cfmVRBbodSZXPLp1kZ/Z7+soU
jvLe7KkkDscrDA5Rb/wen2/g/pfuAw3//JYeizo1ky7cGQYi1uPSU1mGwczFd8iy
C7nMsb1PhBFLgTLiACD0Dv3Ew+hLHHlG+dm5q7RRRrlbTILwvEkUHi6dsHwbvO5A
naxm3cXqwEpITlCanM5rshEtiftACf5lamO8qYkt1P/NHgXjgKNEsbedBvPYsY72
lkwgYm2oh4aogUGOcHBvmGug1aAxyqymRkxbbfezOjn4TgBo7Lvobt/iOpNYz1/x
Pwb03euPM95gQyBHixrxl635yhsaU1+66dfK9O0jqd9y5sxqxmc/g016/jPu/O+8
+TxT614TRY7OFMZDJ7/LlBA6eJ/yTF3OIqfr1LvbfNq2SKoJRBxeHZreekYYvNHA
sP7Gja94MfwtjkdJa4DaHUaX6COgdCZfZjxuQTL8zgxmyke65JZ4Xmfvv1tLpF43
NzNbKvr1PYTqEIeCgEcvadLesMXf5K1UbmCgYy6M3QjsRFUu59abMUmaCQ6YLcoU
4Nry5PHrMz+non2E/Xil5j6h1zhF038TtIsW9q7VLsmDnka2jffvycrtVUywMxwy
3kLIZpoX4nE62U7HohGPDiAS4bRbjsq15ovhS8lt3U+blj2F8XJ6TU00DRQLk+lk
fNF80El1sH7Iacwe8ZZ18K9D/0Uvo9wfutFe3IiVpfI5ODscmARryFJ1EDmE7WXT
aFWOiLvli6FZ0qaUMTMd1PgJH323YOtwXOzp0t0ZOe4u2t56/LLbN2dKNtXQuPlH
8Ha71KKyj6dPlaYeAWeOHkYKYUpsFsZ3b3ntFAkXym+KHXgRuO6Y5nQthkVcqMO+
FU/9+/VrOauZ6Iiq9m60JJOaiyKYey38njaY0C50i+Be+bG6vwgrt9IlWX46XrtU
qW+Mz2fgFX6N4eunEJ7nQxJA0LHeEUu5vrLcxiE5n3mFMuhtTAJ0tvMSfOlJB//W
fG2E1RMZu0Xybwe31PMs25T5M2LYG+O/bXqnJec6AwTiLIOhytMkT8zmr3k7tOrC
PvoIhAXmqucfgu3tF57QSDYHkjmvQY5RFSS/eq8KV6loOJyGrWySMBsqyd5NkyKR
LPShRPHA8+5t3SjJajRXW9Aih5urL5MgGb2DNoJ62uaaHJMKRt/39MtuYIUWAAo2
rXDObxmRtL5zw4RfQePMGgkG1O1cwIZyqezRJuvOQ/Nr9sUTFimUOOVeS3WUtbvq
s5fMk80hdrSwQINfcgGJbiaJAvVT9AiqH59xx/jBaU/OGRkrk3ASCzrORfzzXgHk
MTLRtgu4LJR9iri/L9aTXv6JGChXxzf21580ySXeNRna5uN+vF2BXiiI5x0fBwqd
PAZp5XASCqo6Tc5CGudYO/n9yKwTXeba4siqZ9jry583W5LiY/6mepwoYqkY5esz
hxbw5T97vYacpSbh+z9Q8cgQUrfRNj7kbIQ/16+KhWDgfRq9yHTRykb6DHks0y1H
V8lfmaV5KmV9tEWkbRQLZxP1uDqbtIa1Le0I6b2B/UHHzmBLZ+SLZjWD/wa3ijRI
u+yZtd4dO5go6nDAUKA7xqwGq0zkdyey9LxylMHfMHD/xI53dSBcyebd9C3RUhF0
879RQXR4V6f41eg+3i5QOP47zMezPby6fRnP17b6PkIlGwawCGjUMBDLvF8LoHTX
aQ2T/POfGECuLyctRc3eaKF4i8mjp5ndXrlyh4UVwX+o5+f3W8fub7YwEz71+PdS
bM4klHWkpuPsq0er53Ji72UcjZKvOzSurcIzBWUa5/u19Lh94Saj6B6WHA6FitMa
D+ELTPvCd30whiD29Bhs4QU0GCNDUyApc3d7AWOp7QfKMhO9+Y4TxfDH39nq8tEB
HeQjWVnTzzSY4cC7IQerDD1yRkatMmJNuxmgNrVooSD9apocfVTe9ddmVD3gJGr+
Ch1PB+TsVC8XZVcq/HE4WG/v8jWpECWsYcTmu+/xvZsf0NFYPWYtdIWUUCtuw9p9
ik8MUYHs4F6fGOVY3xIWdjyw2SNYZ1rrj+KGZQ2lh+al69flGwZpFctMaSdLLJSr
ds4liJL7Y5Ai2N2FFEg1K9GE0b94WqFCTVkojXWggjNInecGJ6MhRjmWuPx4i6Na
FcyBX/1Im94EB3SmIefzNnfc1FPtkM3RgRBjwNG1pBX8xHteU8FhuvPn8PVQMfTC
KCiUS93j6+BrPvUyEskvkBd/FD7rN4t7ckeswYuxbJUboNC2VzALEwsPjSrkSAUr
mbdYxGaBu3Y2jxkZSAOSpMrXKIiYZjTWhZz4ByUaJcg64NRhzDLMPKQW4D+Jo9Y+
FziIyqprD/gnaCnJm5bd/oGZSuCX/kLqmEjOXJ3IWjMr6nL8MKar2yOncdjg6dEP
Duxh06wnAJxPyz/XUsMtDwT5ibtpBOW+/mqFpHA5uQ9UkPQ+vyH5hhXRFN4z8AFD
nwQ7x1xQLXaF2BJb+s5xLDUn1RV4WiMmcxlqeJlhAMDHrOeFBDQJd3r+mny4X92Z
nsBVXZsTB9DWHPrUEfYpL0Umu2TlvZX/J1CV3VWDF/oaxN/+0TdsFSDZc5RSmOT2
em6Z9DszuXBtemA22Gin5h8sq/yXVLvfDxstbRqEi7ZBnf/eUsvHBay6EXKY5jlz
iolBKc32r+p08ctm+2IpXa3e/oXJ3kIkvzEzSBeYyOeCMqV5lX62O1P9qZ5sDPRx
vTFJP6M8TVH21TW7LFUWPcodiTQSBnUlT3i9useVTFXj+1ax/hgOAmewYETwiRJg
4ntckHARpv5dLvWnuOlkh4XrizD0rcgEOlTbFjzowdrdadrnmIQW8XyQDDMGkrmV
s1j9Gu0fXZINus/Z2hy+1nFJsqbKXAwUXsiXHrCJtE5PJP2yvClYTF5WarzHfLnG
PrgROxpYgZjW16xy9WU8gygMQKHGqzzwsGVWYFb+9DI19aHrkxLUuzCzVZHBdDM1
eadhMeiWvMwcfDi4k8d9XY6r5QDiuLbFv/kTmVOsPT/RHi+Ojai8+AG8Y8o0RKAb
/H6OGxCURYifwhOEuOIHFkp8BiGDb2bKcLxwYZGk35Rbrh37T43+hNItjoDX9vof
UJUnI/u0tqAzuLbfb3sdZt9s0Vvk5Qyt7q94kJOJxnIntTpGMGICABxT8yuB+fNV
iDia9AqEK+uhs51O6USE3oljQKTuDM83jKjjG9gomzWFxXF4+ziQABjEqZMviZpM
SufS1Bi6UZGfRCVq/xXGYVgUabpbOzw/2VyWz613aHzgZEajgshh7QASJC4187Gk
kXm4Q16qNEg9ijPXHJHzS7XVoKuPy+Ih5/ZUfLURNbG1Beh5iwg1k2vQf3LF/KQE
MFzYCW4WoOYcs/PRGZrRjGtcW7IhMGAkzp0TmlZKSR/BPSfF17s0yh+O0W0Lj+ip
xDnTz4s5e0l4wvGjoeUuiiIMtRZYJXIRzjIKbpFkzzGyOEscYDdS/QXon9z42+3Q
t0r+sH/CDUlYhwJCJX2ao4cw1SugV0u/BlA1Wm9hYS+EHZWeFpJWoo6E/DOmpOMb
xOlyqoqobadT+O2JTHv5NI+4K9JJ3qmxhpJZovjU6aENXQb5D715KbFu4tAZcGbb
tde1j+oAjVP88RIAUK/RD+rfcAPUL6Kmzg95b9aGB4GmR0DxEShKmPFWLuP7Zkli
4tluDhFIDEVqnq/CCoH2gCaQvYMV7T/+cTK5ey+kO+LQmQt/nMACDB7nGEX6pfbp
OLJmHB1Hj+lRxx/m2yRkGtflEBq8VWJ2HRcSbPqH8aMAUNwwHt5Yi5sO56VUaYzs
3XkSxnCfEREA4c4bx0VK6eA7zDYPHr2DN3zBYdTTMPaAyLV9jSnzJuVjCAttZpSo
L9k7WBH+M7EwCz/FmveQZwWadhHtR/FWjQBsdAAdyZ6kqK/KjmkMC0+VSIPtf7dC
D+fiNUuFosRebCpDH7SVq9jsH0BHmmr911Bl5NF6aLtgt2zAQ8tVvdRWaHUqomaH
gLIfV8QRosMUPm6j4IKaDjTAJhPga14osj1mZ1QZ+tBeQjb7vnbBGcVLTCpqT9+g
Z5OBFoJV9x4uLItIC+ILtDzDnxNYal/rTdlXvaBL80WTACIWzixtkZOVftzWkRXF
qwchC0AJwngNPH06FSpBVE0OYt0DZc4SkoHpey4i0hZ9PfsTBqr25bXMJxaW3xq4
51f8Umy+FTSO8U5RpOhJe37jZv2tsbRmzbFEQi+qGSlTb1IYt2+F5yzRtXh1+Y04
NYxIKBa7gIWDNzM8zdTAtPDr6IVfBcJla1jef3ENFXp7J5LMamvEQaI6z0S+RYaS
iHcj71xSjkUOaAxUZ663o06ML/jHV9qwfiUA1TBcvqQnErxC7unYOzHP//y95rX+
yuYdnV5tUPFtiNQ2CAhaGdW3SYvyFM6gcB8ckRLbN3SSMOr8xhz1qEQtS5p21l0R
xWS3ukTGBP7ptSMQh5INH/2IEWYy/fMXB+/Zc8bTrp0HvdqERjBZxgKtUphMesQx
hlx+fO6mHKBsh72RWH9RcBnMYGFGcR8rtIZNdBJozOVs3tYaY4rRviMwlo1L52Sv
rxi/l5jPYFPmH8Q6WOrTB6KGS0NIh27RmhoQwo+yCYlR3beZY79qmq+QJqoZsFi2
osABE3xPXWKzofY6AJQ22mJxzwWVxk/5fb5KZfW3kMX4bwFbI2VY9T76faOOJUpl
ZKohbt/kLFfC/CkN3KNrIP2qXeZ53wMzJG9yvYKCjvo0qI9xixkutSlPuD8LiXYv
h/jDJcBRY6Isf4PVuI3oQG4HO5kjLB3LYbuoCb/ON6KpdtzVU5oowDqLc8rW52KL
p9ixqkdGp9/yp5vRav0cHUkLyHYCzMXmMN15jkHZ6CBuE3clnivzJPM+aemVboRk
6nfvUICPxevtjfBypcG52pbWAVhQDahwZyEuqAzgJCbAS/cB0kvTSYRuwFIxRD6D
JTpJIke8MyFQqiUuFrBsRaPplbcvWxhTE8gJvcWXPHDDL4rPaLmdGHv3+3BzzRtk
+YkZWgRLgdpWdcZR1p7nmgb403mgctZ2DHEmwI7zsAdnY1UYgKEnnrEv+cLA24t5
1jvllgwFkhfupqg6sbEKRwREIPKgwELsiVfZKqVCO9XGeJKfqj8E3L6kcfZlIIOD
o7N3RmwOTsTaiT6yzWLO1laZQwmJ/++rE6h7SwzKcwCgPtZKdf5VtKkc8M8tRZQ2
cA/EjIHpVY0FE6sl+aVwR50kdJAcp3l7XmpJ/26fU+Y96UZ7NiOOLZ5SneLTPmLG
wj418rDXF0o2dLnqi6RxVEemroSjSrgSDpNWrQIPHmsa7lOH3Qhqa5c5e+s511j7
jIZmfv0rox5rM00WOQ+romi1AXwuA93hf0rEDJlMe5WsDl1dFXvuMB1Mird1miuk
SwpC9DUFeIpoG9f2zZycyC9Z0hTPbdeljzbKCJi1yhhGB/a4Q72vJgdYOGQUVdUR
jhQLwBnlTe7nq2QTkDMUbaztgmxzT/3pQiV52RlJ3MU4/tSzE2RGpJwMC6R8ZEoF
mwK7yEU1GWoO/rqizkPwiXkGpLGiy3/usyCLRlRdUdPJCS8XdG3NkKTwEXpG8n54
qPsix5/bCfuc0rulj78EUGHc62z0QLMx9yBtnC8WTQKYA4xKZxDiLfVtFfjKpkev
7uqky04Buc91+FzCJplKRddvT2fngNvMJg9WUEsM/HTo5eSOWtbjAePz3R+BLD8k
SJan7otxG8EHdjg2feoMNKYlzz163wwFpeXcyGcZSgrl5uoqO/QCbHmpdmF5kX3F
2wzdpO2rLj+RoCSLIEsyu0syQO1y7y5UfPn3vQW/3EagoIpa7w1ZFpUVJBxE3vRZ
OCSXrkUHo8+hzvRdZO51o41aIOVaZcragGEPo7f5nODF678mlr41KHDGIxiDDw/N
YQPMtnuz2MNkL+5rkFWElpeLkhpUr+Aq0ZvWSC79OFqPkhAdEZUi9LvBFSjXA58y
23Qc4Hb87G0sxQ7iO/aLa0RzBYdS+Ls/ZmLiBp4I2DfCcuUtkdJHCYAkD+V3muqC
gj/bTbfqv425FU9nqvIN78o5Dr83PvPGmvMRlH0q4VMGUZGvZSIfnzugZ6DPmJ+E
E1GJ/W+8vDxYMtMw2F1q2dIWWGCQkTRw9memlZ/iS403U4tpMJDOhp1PSTDtO4on
0R3eYxOqlXXdh4macJbp+DRO40uZFszrDuBqGRnpU2XghgKAyCZw9stLtV9Z73wH
S3FVxtwg5FPE2a2dsFHMD2H2RI1HqKYyvo1b0u2dreA2S2w5w/xHVNfd1cyPagS5
beW7dtxsedGNu+99e99lCTvBC/wWdrDIWCBirTiBLIjaRKxdDBQJDPIKqpALtz1O
ejPWUJo3itdKoQ8jwEvHuH/sy9Zusn/2L33TpjszeAI1s8OjrEERDJ7M3s0f/NMF
K6jK66G5qL5IBmxcKg2Sai4G+7OUr77/Kz6/uuf+sw0ym4KiHgg0k3jBHMf8rk9r
XVApxIWk/sw24HZZzunrHbjx/m91YCT8HjYLQr9NX5rlaeNa2xkFIzHaTWfBDz/j
fW49agu58P/zAIZHW5GJ1MyyfaPpwhk70tbAiknlgH/moP8GlT1eQ5x2GN8DC5bq
JdjCZwKkLblj7sukEMmaLJhIDAmOQyPSm7n+Cs+5IgFOSm5/VqJTPVIpZLxde6Ep
v6akluMIwmNR7zCfGK+oL/Pc4r6dzqFBi+eQuscxDgBxM3V1Cp0R4GMBJe2g6d9l
xVZ5nKaWP/cSUiN4rIAwMY8HBtAPKUNbaV7RX9AX7bl2JbqfSmv12A+oJ3fPrICD
b4sKAA5Urb/htAE7HkABncI74CX7lpgbENatwal0XDRgLNPNdbU7yGaPe0tVqzmR
vUAN+Hydi6HV7M0mmuvgts0NxLrWsvfvVLif/EO0MOcEYu2ix3WlxF+OgmpzNe/F
/KNaiXIAvYQL7ticEvgRrDHyM/tFA7C+2OE6dpfQc8YdVi/cVIyL5yfOWqij4j0I
SCSVDrX6U1zWU5qqQFK9f94gCWuOxvsaK9KtpZFf2/DmZfVUDI0fJwstRuEJeB13
zKbsubNCSvgLGM0qP7eJYqVUrjrCaJB/s+W0jtMMqhdSmws2LE6GQuXbNl71IFH8
lOChgcLsFPdOovs04tp8/YkjpQqB8Pu9+hbPRoeHnBlbYtAywtRaCCyGcsItf10X
Nq+Y+tG5J9BBxm/djJOQ3eOOWFBzXg1QnIvq04zO+GoPR/q8DUGP8ngHHu0esq91
7qD5mF2K9xek4XDrc0Z/rJwsp+yQLecirfBEhKSnOeWy5z9nClQr+1wE1wrpv0aA
Y82xvmYhVG14saD/CSKSzcPAHrEvK3Nxlv6qTuGH/iwk0zSt6U7Yn4Wutt9uQ6Dl
2bCCKn9BQbsTOEEcNo5/e/d7aWeeVNvcdcKXPh3jkIlrdvul42eCjg2wiRZozBvH
KlrigmyrszMa5ST4DsPDSdbLiOgT+hEftB/aFjcmP3nPQP00WuKt53gmVPbOxw14
wu1oVAMQDqIeJEbCxc8ayFm6+xefRSQG1ZlsozkDtmTcAEXgMswuAmvXcM+mM7yc
oTaNv4yWbQ38FcHp1136HeXtUC+Z0zX+evk1Lt5hmYmFdEUr1k3dg/fTf227dh/3
4tkfVRH08t6xa/qw4XMO5zzN0RpupFp7SjD2Np4nstoqE3riTGvXN0iL9HqpFaNt
uNIlMRnBCi54IXPyJWmIKg8wNNxX2lUY+SbUdMm0FLurhMcNBLVksGUlQIinmQOY
68YDbRM9a1lZ1Ij8n5SsUKeLSB97o5846COjWGltiHOeHZkIjNKh9167xgQ9vfDB
0q2Q5ejJXoyPZYk/zZUj+PUE+XW1+el0afNBpgCwfNq1dN628144O6duKNZtp9lH
vZnyQyImfywfyfeIQFRaRWvilLqnwp4u2MwWysNDaX9+uXtZ030ElUQzmJiDeak/
ZM58UOWAY1xY2nSfyCvuV1fYG/4l4pXpeeSO5OaKUqdpYrorcmd5yoKvWTToeQah
eoVuG2Kmw2HOjN7Rgl4Hr1xm3s4l/krp1JW65yn4rsY4xy7Mtu64jdJaJ4OzeDjV
TSHdIPu7Jw2OKJXmjhB+iiGeUsmvu2FFdEqk60DGCugicU00qlelH2pYVHO5prVj
JaTko+QcjKwLzNPZt12mXHbbcYd+9SKugbtwpOk5Igjgj3Izc8wWgO7/0Nb6iiHp
hxngT6DPaMlXM+r6qvWK5EofVjh0NOkalOHJyDCYQfQhjpLmoMAiJLy8Vn/FYb/P
UGyYfFulBgIochutVkYNGpAONDYkqd8boBVEy7Iomt36IGOKP2ZKO1invjo0lUaz
JPEuPWJB5b1U4YZ2IMjzLicGwI+66nT18A5u9mSPKrpvUZ7SoqzuuUkfKu6dPp7P
tXtaRuBgRg7Doomcy7P4hGgrLcfbhY3uxanMF59nBPRdfE6LMpcQ72M1l0WuAeBk
H/ONRQ18eftdhhZWFI+7oZrDLPB8fcBsQiU/kb+KBI5PRrIpl6IxLCaXWF2WkHOB
+Ji38wblQC2i0M6ajHHQADMi6dRYsL5TkHG85qHXRL6I4SVZEteaZ48Gqx9/m1fD
rn9DHJ4HaxcPNxNaKhG8Zak3RVPSLBzCxXDD02IUThQ1iyBlGQNDxl0Qy068oEk7
eZe8V6jlvQR/N27G8lKrpWmwnsRuCiEfcgZNsGLx04dauD2Gl6hhiYMStvfnDsQ5
dUiXmHFbUesc56K5ZuZd/hQWiSQ2B24oWNnOSfJ776dxuWa4YOfkNXyBKWZ0Pipg
dL9Us/81l4MD0M3f/2ze1dLvj/4CdS1DmDnd6/9v/NxAVeqk9jJtDJT5rHjxidkT
tlVqrwd5XMR4zk/BuJJ0OqlcuOK01CigVdOmLm9/DxntAXnZS86lK2AaSIEhut1A
IYBPQSewK0FaWsXYuUh7hkj9fowxfoEPaHIapj7Q/ZE54IMILTSNIV3/+fXAa6wU
AjIAxCfdj/qXmBB5HKAdxwfqwvQm8x2+1OuyQOB5He3gekrP9IRSYuqEXb+QZYEt
uoGCv5SRYV9Tz7Y7JK56A4dvx4/h6d8UXwVSVh88aYWZYEuplEqy8cgYx1O0OFk1
yfiaDvgi8zGGNcoLdKremgpq/TFRK77wnGmMpNLg9gK4JlCCwL4OLxtMpy60p15G
t7ZBE5yd+eu6YhdJF1/TR7MN44BgcXTBSXb4XK8dfhyKAn6y7DGTy9YdAPCJgnI0
MXtzY0y3iTZdFmB8KAMIn0a3GM7wL/u2SHzrJSo5kAGaP1wYFcMAYg6+mkw+Vfwb
+/+VKBaR/Hrwua3Nit9vLrx1BavFyGS6CCyw5XS09eGtK8Ds3ASN/4Z2914TSgMp
uM7EyH7XinkSzD4BAZd8iKBEThcVdYHUGBiLv2oxEeq9MSulENW5rJaBsiMxv0Gp
W/C39L+3D8ea4BhkKpMY813FjyFGK2m2FQK5pb0UhVl8L1PcvMMotT8WoJhMdvgW
hNUjU4o9Zg8tLD4iPpT/qHRbj4gxXMeBp8kE5pOmnyJsten/vqSAWpem5XKZG5y9
HLsFTJR34JxjH4JMjHuzYqzyvQFFrd5IX/wtgZbRHqMD+m10pfLTlwxnwwVEtBsE
N1CvTxzvYqd66E4Su7qd3BpHZBvH6WuKJbc5RrNP6gu+Af9ItsnJPkUHGKO/A5uj
H99HnIeGuh4f+mk2zfSKbOp0Acb6ENmtZJ/udTD0H8e224Hj06QVxRFdFoz9ScXJ
4ozxQXC9rDLalOFb4mDH4XQXrMK6FfDwarbTOMylrTKGHnMmFV32tyWvAY47R+V0
IJabK3CrY+Ty3rCIlGqpmsC+t5RaNQHhpe8aAJKCPPzHsanxjB7MZDEy8b6vZ71F
yLh9ihHC3P7M7sdTsCdem48jjff/hU7rvnk6DpgtmHL8sgMLl7EXzQP46tx2uIQ1
QhkvvT+mChZpgm5JrcJawFgOIiez+7CsuVLey7TPAMtGZiND7n6fM2nq/EbMb9Lq
N6bDRomoA+WJxD0tl4PAmZiLzs8xgzRtJkAxUiTOzrKRraqO0S8rpY7/vWla7gXJ
DMZlLWosLIXCh7ttGS3Sx1F57/xrjRKkwOIq4a8nI+0QELYVov8dy/yfvddT0L3m
4I1CiFb1xZ/a9d4V+cj6fuvxL+5kLpzR+Ds0ksN5FtslRt+wOziR7cJ7EtHro7nQ
ueSQgjaM1sqWADN7+DAIJEgDgipRrd6DfLfTQ8nAK/NtxEE+9sRbkBhQGoib6pmh
NgoTJpsI84FUxg4sz2dgthHX5oDxVGLGYiAiO2/OwaiDoVpnN5WA8v1wwhLfwViO
MFMoZMUzjuu2SREBVDM44PPmJqzaBsm/QroVJ3FCOBy3yaz5fxOhJBSwkz22SIs6
HK+7ZYgTKw8MIfBOU72InTorKWWnMUuvbKerJFVWjltFs074d/dBK0kwlz1kO/ky
LexKAXw2GbF7//6coejY2NEbeeIKoOOAB+t7Id2wY1gTRmXXnabEJJDtX+EoD/D/
hnWzpfUXgpmBwDICw+jSmGmR37uM8pM6xfTdaci9LzMsqqMw/65HZOkoduUwcipo
rvoetP9D+sPDmYuXzqZ8rk0GG3Yk/S6ZcuNmcBr5exX72dzeJlZNB9BYRTZwYF0+
qeaJxn9HPsrl4DmfIz3Q8G0nE6i55RIoM0rGXcfCtbm8cRvI0BuIvNx3bJMddeK6
4eDjPa0AgTY/bhUYulg4OEBTiPttES/e+pljbSX2hSEVDyAVzVFUCVCSiTmONa+k
xFrsuJA4D12f6lhjtNEZdleNWoQY5V+fjAscK8hJk6Rm9R9T6XOxkAAxRhoT/HTo
kSej2eclmDzlsiHWNmI7WaIv7+0HXNuToJr4dVcFxK2w/8+JG0sHG4vSUaV5r4X+
n8euU7/5/3ij/WkSlVpZsCDho1xbLehY+EnU4RPGwxSRf+RsbWrIZ5yXdesweJrD
QwvVKtFkcEhogaVUKHw+D7UDxDTd3mOGjTl9Qdn/CuXiV/54W9V/trUVEP1+m+MQ
DSRHgPNLiEFOBtrfhhaLoHgfOiOyEzaRilxIP4u38JBR5FM4Iy7gMF3MLUQUndM+
8AbM4gsopsunytuoJ5ipabMFmBZ7cBBDOgKouFZPlbjUSJQ9yopzf/94zi5W4HdP
04WUfJ+yVa7r3Yj/7HXfw5piYMCNwb/vs/6hmDrUZwf8zgcUMzn3zuK9Px2XBYZj
GJwlBe2IgDH9vQArQBS42Agrk212/4v6s870sWKV/IzfZX5ApG/njIFiFXMy2GwF
AvLUXqoutgsHLCfVzUKE3rev9aNB8j0IA5HRUY8KpxBoqJ50VIr+YzpOREN3ERzV
NJAJVrQhMjIBBY2SqwcCqTYc9TImKNNrcLfLjOL6RjsRHgGZrbmEl7oSYJ+hJVwo
SkgtynfacSGMIaO8EPSnJevQO5BLr422DbCM+GTBna6L59LcoMwz3bu9yG/XIgq/
ojYtcGc0XISi1cXvphGY2QTCXnaQDHcsyyh8NhHPVK2bKbbSVuU7aiXzRInsKLLa
/9zFrmmS41wSiSuHd8oTvA2Sc6LyylGHUsf4AuLfpIK1sFlRnk2nNHTNoGL4l6aO
bOx87YcS7deoyhsVGciJxOLdP+EdxT3G4HjOtPd2Spm7SDpYZtjAAjibOXfcCCyP
Wem6Ex7eEP5tNHeFqgn3GP1ekfaX5hnN/tr/YFgUFc7YGP19ZifJu74Oz5EC2ws0
9LyVkJ0vQTXSCkivJ4B/IYvI93YpWv0ZUsiWtTOdcjtETA/YbvPbnquSas8El/EJ
OttLUNOBlZybIIGFzdIJHmjoYeX0UCz6oeLPSI8glXaPqtVgwOpDX9dwaNFt3ETM
Xkj5mMMxQTBpOuqMiQ3ncRkQIzjRmA1l/Gnz2xW3FdY20UGQT9URvmDAMpIyjMOI
a/ji7LVig+PPtgcD3AdoW/uZbk0Tq6GCJDSfS92yeDN0vS3U+GehHFfEdLWfaU2C
KXT99PJYYvpbbqYEpWcnueqtVwJOL4XLYGEg25sVKda3pbZlZd3gzyZv6prmm2GR
OsX+BlHor645OnONmjQU3ZGJ10ZhYUpDljl49v9q4S6lL+J7IlIhB091GWrg5oYJ
t0W127IPtDQY+SFw1z7zZbP8WiXiN8Uo4L+yslaJ5bL4Cra4P/y1l6thcxATDM3T
K8CwmAujCNiCccJIIv6MHXvpZCOr8DP9DG4KocpBWDLN0IOTVyuI1eFDtwCsMo2J
FmW8vIyR8KeDzvx9YyDuaNI0vk4L1svmjIiYngMJKP4HHWUB9s5zUqBbgja5cYRc
Tjj6zcqo9leNWyFgRnkSeG9QhA++n7QRjIPjJwqqWIK5RntGyBRreXhlDrrA22dS
USYLR985mzlj9XXZ7qMr3M10yYKqo0fceNl39yih1hNS8cglaKMI/a8wRSGbnUw8
I7hL/2JuzZ/iiu5/5dB+nri90AccPMp6aeESh83pIfixMVDO3Fpgqz5QWKkKIDA0
s5dfU2DydF/OB8sFF1qqKmJvczbKzhslQY9Hb0YmtxIB02itUW1OIjfZGa5EgWX7
HPEEz/P62hyfDWnHg++/H9ZNi4VyiS13g3fsa5TME63RoZXGoCtGaGXRpvTqU6sR
2DjNDqpMjWDRW2RBprINvgEx2/NYBpJ5BkXi7Dh1OMs=
`pragma protect end_protected
