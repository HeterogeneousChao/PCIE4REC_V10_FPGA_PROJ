// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:17 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qMs5BEPHmpoK7Bxl7bQZ9woawTtefVApffm1/F3XlP58XaJiyUTe4kYdRmRSmLGt
30R22ch9u/1NgnEotyetTUdVrRLkkM97X3OBM6CrbNzTWCu0dDpL0vjGb69cS3dr
Tngrfn2HZzedoD/T84kFQ5JK2Zv5Bw7qIcQFYftVDDw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
2ejU8QIOULwDB7R/1mgZNazcCptFTF1MccRnAv+D1j2laoI25z/KJH5ZpelZbEbv
AG4zXvXfOwBWJ6AMHWuYFdVZZhtCw7itgyie06Q0b1OcXUzmJ8bfd9Zu3ETEOdVo
m3YCTfAJ4F4Yysfdj2+8uYu3kozfkLG5d4Z2YQLW4kv/mQnfMXgEgVGUEmhyJ+k9
M1bIvQY2W7e0CQGIk/ppXbaga12TPajyfBI9J1wylEhsAwOEOXLbB6Ke6UTxz/4G
rM8JOu4gO6mqBXE9u/PMPMwK9X5cpz0Bqlu10aXFFA9T/u2BMCT4QONyVdNZeTBU
UxQVUs1DHSxGn6KnGLX/WeVnTrcRnhFMZKGf0gQAq0bJN14RTLFnpM9sJh8W+Nmk
Pgyi8VkKiS7/SW46+99MiGE3ppezusj8dnd5PEMCGxf0DtzUE4EgaqUZ6A5MTDPq
DEQt94LFoTEAkjUiBv1tFdxz0YeWN1qQXMTY4xGZUyhH77bMEJb/qyJKS7H+Ficc
CXssJzXcZxpWTOY7u8UYh5oR/HcIoWetUs5Ybv5CiRota6GaOtFxmGUWU4nXvy6A
XByASLuwByHiE48/A4o8JP7c/k2CF7K4+N2fkUNV4qHfgmomKV2gdCFGuaVi8w1s
VpO8RLyfarOuE0WSK4v10kwsqaf31q+X+uLGb+RJ8ALIdC1YRiP+u8sJD/SLY/iy
QSuoPnHHr80+bcoQv/LvhuLywz2erm+U8VHDUpgCxqIp+34TovE+O5TVBRWPJsh5
czCxfunO6irGzGf4Oh3b3yVp5pNZogM1rMJXOd/frvCfoBSp4uR+mkf0GKP6pf0+
BpFUpkbrGwLs+dx7ndAhBUCHukIDi1eMu4S2Vr4uI/i+Ha9sxq77cxMNq5TahGcx
n4cYP3zzm9JhA5tDnQskrAegaGZ0StGInX0gIIhy1KOWGOpY+jXDcxAckJwSzJTC
9rbwT9BvOle3PPHxM5W085HguLXd4mINfFlDxVjjD6UblNcBuEbw1SZCD76ZASLH
TQsc0ErRybzh7wLWthxxrL2XN5RdH/wSl8c+OEDLrvUg0hWEQQuhWe2QTPxs9y5O
gYcostqSLa5dcYqSBzUnJUxo20ow12WPAGyS1RvcpXie+PYDUZgR8JkSMuz9SIWm
QR8lPSfjV63eMEqOzNp+b2KyipxEkrcPNGWBNcr6SVRsoMYaBQktzA2tgCB9tca3
X8d+cfhFpQCFXBKtNJnDlVSIgVr82h59hWSFI8YhEYRcZCvg4WaVWTzfx07NOq2M
i+kEabctJbyRLJjmCIHYozmRe2MmIX6uFwFp/uQNnY4v81U7pXDGmMgO+XTsUrbt
K3yjm2wuVQAw9MUmXxPxM3DteoQ2nQiDycvQp2kmabq29PYbVM6KeVx1nsbDmFp8
wdyS75TbU6TKrxzrnHovOpAZ02RI8IqaRoSSXzyB7St/6LL3uAkzGrH/nOuPvMMJ
4t38eY62+wPtCxRmlDmBFVyCrcwZR0tq73Fgt530wRwhSGvvNxhkmFjyaXbJ+lHy
tlVAqLwru2HBm/lG5lQNHZoIlDw2UrEPBgoQKTDCdS0w5huNHHrp938XucDxZbah
ZxkPS8nMZu/OlMl+Z+nvmnt5N9cYnbDkct8jb1hHOsKQ7TsBg1GTvALbBLlJ+ibd
d7KiAzlZzH3a+06tKuKmjgVHc+p9Agfn+CH7rgtsbWUgLbjI7XzT3Lo6v2sAiEsu
hdp/4X3dXZNbD9O0xGK4+FxzuJgrP4Shg7r+S3moPLbW8mtf69QQUoj7vSkoUyDm
IfccRlACao0qSMATFRBRnKSeKXZUhUFkbFJkVMgR/ZPFfLdJcHsR4gVYYJJPwVb5
2JnN8abizc8envLZnwDdGn3gcifv5R+LO+qcSdgmdfq15wDRFtHRboL4zK+CXi71
VfjAHoiPsby24OQUEGPp/enGlZb2zrmeH0AQKrjwoDBtMj5IbCNr2F9CQ7RbnBvK
S2iPcae343skN1tDWkyTtUF8EDzf1M0KzsujpAmjJ0SBY356pSiRwNXdv/A68N7U
zmkWZkJsBtfaX1yedyOPYVpGekI6By17UNnaUvzsUQYdmp2OJfT2fYuLQrgzn805
L/u4VC5RsYGA29uCmQBhVFuwJhdpgyWnUynpT4+xw4gTuqNwHk5hEot0KtccD+a5
i44QTej3np0hZGV+aBaBW7pgLAwbsdf4P6UJcn/v3Y5rwWc0lhv0L8ONTrB1L8yG
wJe8rZ60973n4b9Ma4mW3KG9EjyYsVWbsuwSvf8Cb2qhjfFCJTvhJCiA1kCfm1fQ
CgZ4iiYiIDnmUIBsOMyxBJ7t6M203vxabBydTX/RvQTrve/32auRG0OdTFTeBvQq
hov1fjDI0WxTPxUEfvMoCL8B3zZ4gZHLA1j2EUxn2fSELhdNeXBxIfpwvlq62Coc
CoYUz3Y8IdHy/QxJQeBFqwBeQxeXwPlCjwKtsKtgzwyYFBbTws1AfMsN3sN6Op2P
sXDfNNOhTEusEEVnZDe4Hh9MJ9/Xe++imdFKDl6Dc722zBObGD+wZbN67e4ZivXt
VICNF9nYv3ax6fL2lQFmxaiyCiGlp942rlxNGX+t3DmVZqVQ9UEVBHVd0uPHSZo7
hb0hbasJtb6j2R+8vrD1xiJEMRcbzmwW7QxxlAwQ+YK1fg3pzhoEgXsJudWWHZGC
osCrIOzUpvJukiAvOcIUTK9esstmbHlmSHcPq8FDxtIz0Wbmv15z44ydxH2dDHOK
/R05dKdug/1wi18ZkaUJkkdB2Pxz8ZItILuNf8adbZX36P6JaZxIYpuzMNypnBu7
uUH02QjTMtYUm3QYQE2jtKd4B03sevlswX8NwLsh1OxvI6UuE4/o/3Tr0d7RNoFi
M67+S3fUYuaFVJsM5r3j5yAS509aDTHhA8aii0CSB6GOJPf8Y/Zblk0/y7NX3Pek
MZ4nGoSreIF0H3hlTEjpdNxQkLoiheb399BFWjb3z0gOzzEkwp9XfPYmIHk5u1cM
C5G3zojEsaTkbYDljlNuaFuyAOjHVmAVsWdEOK9d46zMh5Pr0a8n1KPByOSd0tXH
k6/AGakg9nAwlqx/STEqS+S1XgNsho9mi6XvugfayW1h7JlYEhRrlkQ4Lg8BtapQ
oi8xL/SPqZbYlSKQ5FbO33zRRCT9gZM0NgwzajwTso1ge20vuDelxVfZLQwtuOV+
A8pysVqJVHmHGq+tJlcgwTwrPq8Lzf5qWH6UFmG6qrGR0Xa7JzK/g5OinFG5Wa8G
ug+NOyKDlr++BJ/5k0DroC6Mu4/Xtn45jLL5DHyqA7rnaElT7C5PKmaC7l3F7mSq
20u3BEgZkEvK7FjC1afMyQEKZZfYQHO0TJ/lMXLt3SPfG3ufmyv8NN7NWvM+WTIG
q7gcwmrm/SU6d3cKzJVjVlHdkXmTEEGG1Aw6XZTszV/NZ518Li5QTRWkAjtPZazc
eENc8itbf70+TT+Auw7YBLpJIFDj1/thPGkzbeMx6kD0ZhuCnYmEArxQws7ovvru
J3DCA90+NgY/5YqlLsK0f/iLyM2De0gxgksnGP2ypLduXfd5Mcwkm02oyR+80e4o
6dRkGoDJpAu+DZVpyxG1eLp8YcOqPzMQacsT2JbfwdpWJErjatodBXPJ1+V4vK5j
ziwtvvu5jOdRJQVCGhcmgTkEfCOj3kU5zCstaEEqoyJSHUOsgm3ssuGMJFs22dyM
HHWhMShKXhIUfxveTCT/e4auyFrHjWfTyo8ZzuxLNYuGrLY+MOaMK3tbn/GimNg1
LwqZRnH4uxczcyvsz1MJRtU0wtvS3I8vGRVQ4nxQIQiDBDkIB9XWIXfPjyxzJJwi
TRaX6/1x9q5nG0RMvx8nvP6azsH+VCXE3QXlM3Ulgkpu7/sJKzoW6DT/8l38VDcH
9Bumf3C5nOWUy7IRKiFk73czgCsibFypD9+qxUP5laHnQ9z7GzidGtIDoRESKMSv
yBWK3l9ERQ2uNerG813iPkY+1p48tjPg6PZAhfEi7prUkVUOCJV6fq5nNB6JRYre
n0uZOrsfUCEpRDm91nByrnvXVFhHEKzk6GaAslaDzFwGW9cIUg9Pgx0HXlWGT70U
2KN3scvSLgwjTqdU7KXdD8elTumKz+pUbQZhZlFdZ6jDN2fPPHKz2gO4mcKF8HTb
tmUuvIcDzaZUWKVUl3nueFBX8JcOPWqTYxO76E2OKIcjao1C2CRWwNoxIhPrr0Na
hyqZEomaTIcjszMBj805/l/CtYou95gkN0CKHbC6PpeXcTyQQehbqo2ODCwKb9yt
AnSzQc+101pHRwLL2MJm5o/9nCzC2zPzefh4rKPP8Lnno9zIba+BV8bBtnl7EoKH
jv27ThDXs20P7UP/b1LO/Leouil+26LZwB0c1xKi0HLl/6fBnzuFdOpSlDNnBdME
jOsS1xQyAGdq6Yz1fV3+dyMJ4pFHGFwtu5NLWxotvquHgI+BmOigF1xLpH6Dzkmd
uOyDszfWpdjs6kgEKocf/d+uh29/Z0MOqY2Dp+q0cYXyt5PhYPEKwlJokyx0wicJ
XmN1Gjl4VIi5yV7o1BSxlz0NqtFW5vmXmV71L8W9Q9ZVJis+MxKzMvjd+0oaf80A
OT7q/E3eeBUy5YBoN/Ny/CZ8xUDh1rCGeGhOc2yJDg9uCJH4R2wvitWXHe9wpiQA
5znqyIB080dw6SNKk+LM8KybsCEvbuBzRkXuwMHNBXgJkkxkQQJzOGKUNZCmNpUZ
eyHPVainu7ryBLelPPfyehyV7NiuA2qFUMhjIwqzacGt/Afclz6Hzsg4WMRUjQK+
5jdjCek9nQyVTx4aTXFIb7CM6sFRGxXZjNWLRpkns977UnsdgI8P61kNrdZjOyc/
RaRVM57kCQ9BgnxnDkVGRjmpXS1Wd3AD0tnduKlFtZjQr4UOi8cXpsF5cWOgDz8i
wRoUXuT4MpgL+XNaaZxvJedyEVJupN8lryqIch1fGQHSFPe39Enr9GumkIvK6Qmk
oxXiR0PhBuYtzFASvx/DyzPUoECsAbhU8F7rVxAjUGMvLlFyWGmJGMOYQMMsePYu
woBRaMgl9BocmBJDbcDNsI0rE/VwPaaCa6kJYHYXkp0aYc2EUPLQXH/U/DsOJ9rL
G/YR3xgEF6BvB3nnFqUC6TWKTqCpCg8vz0rLKEfKZ7hkum6GVa23zyhBQOMQpbiu
fpvom2jitKG2IcMuaoJHhCul61+OdRGKredePBubBcHbyvrWXnz1qx6FYHryRqS3
KtLk13yVW5FP/Xdl+tcRVdCENK5rNF5E99yTZtaJkprmqHhdFO8G9JH62cwo6zB5
3wwIVsTWvMRMp1EQsoBI3TvYA5P5hd7020shzRhX+mtnwLZOtuGViYTsBH8QgR0E
TAk1wSdPzOsDV3jSP4YJTbuWO9hO19JRzIlWf87p6ZsRNI1R3RliOKXWq4+buU7y
ANkfkA31ZMBqeOmKeJ1k7hpwn2y6sEpg83M1Q55HGRjd7FVxjC6UB3ExlUDL7sjk
szWbmACWe3sJtASliBktvkeEahva0n8c0R3trnmbalfY2GUVTpf4LRaItuKKYQjm
ROmOL5veu2Q6OSoEzsKFE5V0mi08+tomypdCNFbqsfDd+HWwkxx44TbDKh+5WDgO
5wZEBpyN1+cJH2UgEiD1faxqyu0Y9CPmig3GpXWpR2yZbCDXzIv8ijRk8mVB+DWf
2fz2f1wExRGkRysEnL2V2wEO1h9JJ6+ve3domfy73cR+fsRyzlmVTVBd6pGYBe65
ueNe8VV1RM0UgTJLUPHj5D9eNGag/TW3GdDDfp1zP+wifOZp9HZAPz7/z+fFPrNX
h1nfimAx8Z9eFao6zhdbBKW91BSotO0Ktth8bP2Xn2pNJw0sF4hLOPeL3Z9gO4n0
2quQLDw0b7rvCVDrqkH0BHamphWY+LiAaOJsaDMW4pglzrtzxeYnInWdk2DD0c6J
JwVJtp9pdXFo7iUNc/A86YNjHcf79YIc4HfNxG9dChw/YJfae/5etNkaxZiS35XE
XA9bDR4gTFYZtzk0I8og+g2nRdufudAM4iWdoksODDDHYrqNiP4hf7w+dlIFIVqW
SlxnIgAVqnqEk7eQL1EtPBYb1gx97/zAY+MTgE4B4iiOOMdhwWFTmHbnM68GG4Vz
xF5lHmraRkXUod6FnovaoGJpUALqZj3NPi3/4HE0vzi4gsryjkYH0pewIW0GJ8bE
sfM5ItnssiS3MSaT3fGD4onIYxKL6jy5K2erSJn1alnQExmYi/IT6tYgjFRKFw9s
TY7cEx66RMKE2zkf3BkF70fthbmJ41B3AcEKWnCDdJfuNpQ2wdOb8XSHbslc6jQP
QVXD0XP54FqawoDZEmKn0kSXef9mD9JagWhQHRscFqpigwv2coQmNC5DZsV3JQh9
W9AP5Zi95Yqtco3A4LjusoQP3MpEcSMfQKnQrTK5sFamYL8jev0/rCeQLVfblPg2
8ZYI0oZCI/WGHYLDn0TluP/FFN14lGvpuAIH1mIaQsamR+tN2vefrg/2qtsG5pA4
FLsm1+Mcn5cPpXwjV4QNTL3vThD1N5Ta3741QHZIkBpZcHDnDu/Lh+FOfkiwew1E
DRuNMNimZYVTBBBKPHmFEhes4x7x1dzpsUwTqE0ZduM/lbdKQIVVEL+LS7rT5qgn
1tx4Vo1ikQ3yNE8VnXB6Iw0PONeCOkRQPF+aMU57MHIogY6GunJQolcq0jA1kBYx
xnTcFYoDdjy977Aufw7TGKPXz5nVnDBjEdpKh86NoT1JdeziO8oNFAVyu67al/Nd
5c+imyePgvZGM4Gq6er7Yu4HQebqiPwCZFzjbrvetSaJQNDdRZvvic5NeElqt2lq
VUSViPmV8SK0MmzwK7IGPQ3bRbouq5sgvKyPFiqnhjvQQ9lYpZkP4w9W+2IyP8B1
VZHHIJRAryEtcdqwr7HSC3dhrrp4cjsmaNtFDNU1aRJmrLbTA59JrTfru0rKK/1b
nc6pirjkqCWVkeh5i7TQwEnNcogA2uTBBretNcMAq5MkTQzKeSvmBRM07zNVA1kS
BQGgtJrl0zzAnOdUBRTyWgLT6VMOcivYCLYZ1sXwQjzQzVz7J1k2/CS2hS1wchQu
GQbDEZnQfInex9N3yGuXYXtT0ew8V9ZE7Kn3SkvZye/qWADgACMC89yj+8s9b4ZN
fJrkF4xeYrJlu3r+BTcw/OoPNxAqtis+ftfOjMpsprziM7bry2YWFm78PIcDgWpg
vASMBr2nLVjhlg8YcocLbX+v7UP15yObZfWQ76i8KSmA3D3y9Dz+tBjyzBxGXHo4
v3/kMFqIaZXckeMVgvEVoB7yRdLJyXJE8rRfHd+kKQRpXB5On+Ve6g9ddWvPP8nj
naGh7J0JY+GeOd+50lJy9t9iGTsG367ADZstZKTB7ZvROrsLZvIz6hZlirs468nI
tf8B+1t3rUyxcm/tJqeNpIgetGbU7CPnb9bO8XoIveyVOODkw/CYoWQFaxqh0Ihh
jfn7MDdfqWLmD0QHKiWNnJcmFZ9MTJqXTOcBrXSD1a7Tgb62GNy2dYKQ7ZKuyNHQ
yrNisqsZhsj6ztTtZU+gsggTWPA9NTNdquV43sy/1P2t3x7NnVrvozOj4Qe3N52S
HCpYMxsmxtl/tSh660qVD75c2VtqRLrtRBZbNY5wxkGZurMLZpeMFNWRz16ZugHg
vpgEoTlfok7lChcDM5Dvjg7pdAZ1QwtoyyhGdplGmjyFkaACk5Ch2QFT7e7MM36r
RHz1aI/ex/lkfcWbiEu3vGxZFmqXmiPFGLiz6quzWALRhTicCuQG2ph53GACE/7B
zRjVNSE0GXvGRSKObY0IJJE/390f3c8XhZ/UgQji08fmOUVqYujRhe7HIo67WCoR
Hhy68t2o6713zCEp85fxRr96F7mUNkuvOYjSHgsgPq0k5E1t/6kjH0hpm4cjexFa
vvFoZJjl/WNLf1tO67h17/L63r26vWfsbyUVzOLuM/41Kdgyp0bXPjG7mqTq4/OU
rh1syCkgglQH9abJS/TJ/gG2/o1AGh6jPxC87YtE68og1oni9+Lko5QGXnxHYELU
xEj5vzqfukzhkEWsHZ3TtTi2SsQpquL5vAyPaF/tK6kmVJPZoh+HdiAclY4qhNq/
bPuInnN23fanBsC0m3TpkruPLhf8ygMzyLInu0RE71V0+/WKc44wh16FGOPCh/bP
ijgR6YlNGwPvcRwPQ+3glB/4SNur/UztBgreMzJAEQEbmC8nwm2F803O+NSO7qvm
Sas44Bz99TBuFIZ6ZVDj5lGif6q/cWPXtB7m0eyt1dXLJnpjhbmhsI/bzHsZKEzU
MVS3PicfEodfgc4JtFpaLbJRHSsrMM8V+t+UZPpqbWpIJV5dBrk2dgqroBH25XZi
ToZd8ISGFIBrfrzaN/cc7IQDRppgrQKc8ppJrHzbPRte7VrZCLeTUEHaaK1ciGTP
Zk2JgKXhJd7cGYn0B68yKyL5LzXsmVGMNLlse0NcOnVZgdn6hkBgRHKE6YLPJls4
BWNxWs4rMik532OFwdXDq/kPvqlbiadYE4qAQd1ndR7NpraQNwz5gisEDcvEXg+B
8e+y+xltCaLF9suut53NB0a012ffUAg/J/hlRnWJVxKCd6kv+I2ve4OqNvLkvXhb
nPYW+M8MwNBEg9PDnrNC68Br+eVsu9hnyi8toAHW5PnQZD+JiEiAOInK36ruOaKN
qYVQ3pcUlVegcsUG4QA7KhFCj/vK12tc4FpIrnbchEfF4Ay23YcyncyqUbkytDSA
4JC6wWoIn67yoa/B/3LItod2i8CKphJVqVWy24nIqLeAfdDyBxBpMAr3Y1mXKolS
n9AJBCzSK9yibRfxN4Y6WuEbPKOCxeEUtFXtN4NRorYF8uDjINqcrNfipS5QBYUi
uUNAS5RDn99GAiBn1uDJNoRApH6fT3Ve4GZcveyVXVjdqgcbe3IBPLyLH3GfP26E
dBWw042/omvEPSUbYTSug6pHyfqeIx+ewl2hTOIHw8ZvGJmFZ1IYwFkCc3iGFHl1
PXbF/WcySkgQrmEVIG3oFdXO+4NYsFm76aiV/tQoH2AN2v09ojnw/8TRTIQgcG7P
+Jiqbwlh3OBxoziLSE2z4lyPlMxIXbemnSCtW7dMU9gzwDtYAClN9kMh4glokEep
h84T4c3m0ZTeWMTDn0HjE3Krau5tsqD4Q456ETugNPZeHf08Bsa/Etj9J525vBSY
oWO0O4o1qj8FyfVZBtT5ilmocGz/+R3SC6tbOfikbo6wzgPqRNbtpfvRSf6pAvG0
WT8tKjkcCspmaIc2azeJtx1E6f3SsGLlgYJtt4cqcpubrEIYnj9THCGvisUMcYsc
fb93qvNwJyeu/oCDfDZHaY8t9wwXBk1lcHW5evPOtNhlIVBu1xIFCAFhSvZyVHt4
MW0tDvBPNvRpJg9XxQJLDad/jESaNBI7CuCgOuMtsoWHCKPC5CiHWXuICwMOjx5B
hGtDOMzhshZQ07KSjL5QBrwAfrCHebJ3ksQPm77K5J6KZrqF0QOkSvdB3noVSozU
dN/bg+mJv4LKDqOcNOYJrVjRcYbAym2YNplbKZPI5sZnQaEf3zNLsu1e0OAUGdpj
qzCO5E5iyX1fJw2xxFiFvh2fpZng79FP60IjUdNxCQABKWrDgDfBA6Rm79SY5/p4
I79DF+EGsv3To9T4Gpm9Txhj0atgs66wRNGVMt++HnWtPDrlJnvWMvFbJCN7wQpH
LbUz61NgGVLvaWnyKiqWCDc15zHJRXg0JoRwo/FpJve9m8EB4jVQ8RDXS0xZmv2I
fZE7KiO8HQSc403zOpUR/SQcTr774+b71NQ2QsacLxZibFBJDDIa/ZpGu5IVcr01
eKrcsZSBsQ+xaJNtrdzdsZLJMM9Uev4e/94uvjpdZ2wcuLUtUmBk+eVSVjIomOBV
tJyb8bMS74Gn5Zfng2wfHQs7obPgoP88nx2v1Wy4nb/E4oZP8HuSr/whjdzjMtOs
wHIRyuY+6G72AY4afc7RN7GYj+kan0LiOnrE9FQ0x4VfCiy+qvfTtkV+EXmPmPrd
9fhH4bg87VFkd6lmDL4eL6+YHxfn1XowbNr9pJ/CTC6tz0xr/hJvJLCYUjhox36+
ab22g/N1+Dr7JlGyezpRRoqd8aCbGmkRzB7dvKaLnEcxeDPT+Tus9gU/2qcxURzp
+U6aac4FjX6OvV8iygXVDFcmLwLZAtkrCI+HpRy5jg+zva2NuIlrjOAtAYvsjG/K
Zkl97ZvrcEVgephzZhWvAztMUicqWvmNfRaV591SWgwUNm29IBE3FxHtxKcqX8ev
dd/YkyHN6HFeRUsnQEH4enLk8g3SJP3jerOwUkUaMG5LzbopbffLes25ybkc7V4I
6JD5f6foIKwvXeu/3oA3mvPH1eUffgjlMfeO3YQcY+5KH2kfw24KKmCRyPTXju8L
x5EuWwliVS4PmkQa3eo5UoOBqa52Ka7C9MrjHprKqMKYmdQmvvbI8Klo+T7ZUuPy
VEx4zx/9GsCGnXu+B9WdNLHbMWTiRK3SMRUctjivNoufehdQE3OJ2KqmNiv6jZ1B
WYzzK0MX/T7HoFV+UCjA3TQsD2u3g0Y06pWSHDiJQ4zWob+9o/n8rv8+0ILAihuw
lSQc2hCQoZSaGYIeuH7Zq7TWpFIhdgvQBmWd2H72ADITJ85eV+psJUd8r4TmLmWl
j/3Zpm+erKMTEgF2HXmimgPwKncRfW3sCdkhn0W5vC/p/aXUMDxdqcMVDhUkCCCl
rU+1JD95M7ht6jmI4QDR9jbEeLr+Lunnu+puDzJ/5NRWlZyyLgRNMs7QsKnSMrJ8
X5rgBDq7tyAsTCXRWUTCVgDctWh1/lk11ICRMpYnkFig+I1Pr3P57k+kLe4VYtfE
qaVejT/vQr8YbFwUighds0sYe5jX9/4ha0Gz4lvjcwTjOUnj4Sn86KIW3GNISncB
c2wNgjdRw9+gKkMi1J/GeOQ8STZSoq8n7lpSu20d/n5tmCfolFGMAay7v86znILj
W2McWE9ScdLOfZ0lbI5UOzCW1U5YqQL1mMa/j0LCyi3smvG9tthDyyF8xYK3fJbi
eUTSMxGqMo7tEEpjkwAPGc1rjNaw+MtCPkUAz2eOlsjk83+5ldAgpx9oNU+rQ1xv
MY5hQrV5Wk5nCnsvaM3/TxnwYsoeeu9XC58Gezc1FA8iPYVFOEH6QTPeFDMm+Kgw
3ROooMqjCHc8JkU/l5KPGbvstQeBjqaZZlWUQkYCyu/XweSp8io2R2eCc2VL3OLB
9yxsEo1yXhH5QACEqCsL4WRMROTlA0IV1/CO3f5ZV9zT+IIYLNeZUiiGZyZ+HzPu
zfxS369pFtTacSd3K0NTE9/tvFwZTDFbp8ai20l+UcmZ3C+gy27eZRHeTxJOAX7F
SNsg6185KexhgwNw1F2qUuk6O/y4I/pHCiQMq1UgnCnhhJnDOsWFbvnjZ6WMEKoM
LRm+RuFNKSxuDxCZX5x0P5pgpFAYJ42nL5HQ5YuvCVF7Jms/nzEa3awXZmCBki/l
8Q9vJJ2QivBPYRzp1LmwRc0Ldeidk9CL1EjfH6jFs5OlWZfH9k1mklDNwTOto5cP
sEPt4pBfsOEoFCbN2IRGM5iY9GOlthQoZUTW+XjdLO+kHRmtf1HhqD5Ko94HXLia
+B5oSFqMTUxQQP3fTfhD3gIcT+Kh8C2Imyz517XrTBviK4Y7kRnXgwSEAo8HxLdU
EHJOHpxWEO7RvmMAFkuySwlizcjZleAHGnF0hSjLYMiAKavRyihviOjBnvlrcy0Z
gwA/sYOrh7coXuur4bLXhi2etVLQKHWw67/uTih8O2klC1KhsMuKASee9lm0AEM7
8C90Il0Vyvykx1LcWAkG0T5whkl1i1tIAhDqcrzDPkn96dYIoukM3LBGLIOMHvjr
RU+zTBKK2kfHjZmnIsJUiH+p6/LVIZqBJF4xmIx7gSpmhsayGdvAFvoDwTMRF73y
vgxVII0o1oXi6pBx+BrtySgUqnUZthvFO4X45ctbLo2q1LauFU364s+PJdeRWOIZ
VcJ1jduci4sEnPBZQFuD4jLjs6Ej2xSET4sEjYhq26dMSCFWDpBBO9hNZPGgR2B/
VvRz98idUGNpakWBUy1p/teWqVk4GjrBi80GIIVaMT8SwTrRTgBb+8wzBRnt0snm
CYSnn/YZI0RY3JjrCEzLk6eldltSDWGf+4r6Ipg2DuzKSAotLvduEtDw4jJ/zxq3
qczcqyir7qdHntdAGwnjvO8SDjKKEVANeIi8AOPELYjsKq4j3eYmb8tAiDNDx4RL
NywHwLBsQ9FsoJFCDZ0kBkdEEMWXO+9m7gasQbHCk3RQVMxXI5XDMaKVjfVbXGH4
FSkhi2XelmO1ITyol5GSkLlV3gkb0AkTObVrwobtMzfS/F9AeIUJcXaJzNR43nlE
7ePsJm3Uf0dDxQUyXG1a1TaMf4Rn0dLCsPawg2sPW6C90VjkgFNAGrZAlf3bmkxb
lqHNZZnJKivr6k+NjAkFnP7hv5R3XeofgYPTtTZYRKXebJIXXqU22y4Y3G8wgkIU
jgZKI/xIM/SdrDMcv207SfGpBKPyIY4LbDzU/pJC66pEJCCFSWm0rGTn3Fnw1mJg
Vl+Q+gOKGDQV0ag6Ytvc+KZAChQ+jfwYqGiMvkXUHbBv/RI5c3hmULPSn69fw9fo
SZGh/xYYkVm0xjWUnwDxsolTvO8ISfBhoVnLuzgcUsscPVb4/YPa1NK8IqvBKWnI
WAk6l97udK6uSaQ0QYCL6bXPv9K16LMBKGmn269F0Li6swOQ6w7UntRni0XINrbx
xirpxyptKzX3WeooKdmbjt1Qw03DkbKmr05qlmt9L9tr4MKydkrppXE2mtr0opoA
J7UBxKvrNDkNby+RiIxIM0t+R+/XCiU5TzS30EGI9D84sX0sGJ2rGUGzqXd4Lu3+
Lw6kMAy5h7gmPzJVbCD3pZYCrfQ3+JNE1DPhnLzPWvBACf3O93BKTZwAb7Qq2vNo
7gLvlxykUWA7Wm+Jshc2OUN1DxuY6s+7xVQP1dRBOiWOb9ZEfUzZQW7Uv6SRQC4R
yW1Gd8TRuX/pFqNMmasTxqQE4sU7I5sNwHGrwUv5yTAEd8Ejhcnbv5sgHRNCFtJh
cfPpR1tsAotuJmbjm3Gjoyi6gd7FIPI3KzX6LE087NVHuDjqecZ6zkO/+zDOMh2r
sd7rfheFUYIkp3Z6Mu388GJVIKnKgy70ghpxNCS4FrGikSdO7E0WuU1JpD9jjRek
h1yHKVSzhoiEgnJNFYrBs9CXB5DGrrP8wv2KCuAQMTqYeVur7qnVXel/n4JhOXqE
TLA16cYJJ/Z8RjQhF2eSo/cIbMtfXX2Su/6Y0R7McZg8IpGW+i012JivJwFQCn4T
iYjA+u0ythjzOVUvcQY1V1PYCdjQZo38f4+eo3lLgv+ZaH2JV9HtNGK/qWU5Zddf
XinBzPmTcTDJxQF8pEkIDUtv0h+qigTcfwopsO1oVUK4a4nqctDWhkMW+bDwOFQc
q3j5gKguNzgp0fOyCibcXZb3kUIzZ4SsV3hB9xQBt4HsKAbVdCmByKqNSjMGp2Yh
cWXa4hJ1jdE3dm6ujoe8f/A9HGy2O3JCB/xZOSYPeEC4YJWarPnCk3JcNt0yFaei
O0UyFaQiw7IDEYomfx2+GikTTMPxPSIUhy+OBLSQrHqXb735mzxfrIkpf/Z9FCsh
F6NnMEgHSuzDKVO2jhg2/rlGQGcK7XSl96ZLVZteD1Jb08DzElOETBfJGf8cIG9q
oE30LuoDKSK7JmhFogIellRKxuNA7v+3rRLE8MwEEVpiJA3pSRMb2xzNjxXsq8+O
HYCwMYfzQ78PhH3D0bkmwAdzS4L/n16hbpcMSUD+Xy/zJFYMGqu77Tt+GNvYM9yh
7ISsPDOBtJ4NnO7eFYyJZiOfk741xXyvadW12hyBkIwNqJe4Yej9lQOk8KFkZFLU
ZtaGkknY6vDmOywS9j3x5bYgQvcOgeF2LnM+DdNyrbti6Ny0HU1Gkip1JQlHF8/e
KdvyxogK1DTnnnpsxhPTCq3DeiqAR2D4ReX+mtO1w5d3eLYgkI86+79EpHfBfIMh
qSenDvPRrbgU865/NvReci+ohR4KWGogt8zEydveB4X+nXjsdiSXLfwJTDaJvnK5
IY6K8LSHp7psye8dagQouozS/id+s5Tci3jlHiA6djByshTaO8ZdGiJiC311TDar
aOmhvEZ6jWGV4SjdliMnMULHdsHAB30fjKt9V4tQgg/zB2L1riHeoZcAUzy90Sqz
z6ZqbAT6pYWObOfDQ/CEiYR8D490VCmesWyges1kl5FDFqQaUGGOcl3ZVHZwP46t
r+zaA+RTaDB3i1wWb4N+10I1wXsiiTvEuVVwhK70nodSHu2AAYlGQImLi/gdGa4+
85+dGjXNlj8Y0MzNA4pkOtaznmbDBm9NkjwRqCsZxILSEtOAQU03GsxGJ90/8yKo
mjYfBkNsRZYGnemgHXZiu52+SP3ubxHdmyUQPRYpqF8WYEq9XxCQSPaiSwwOPkQC
VCPE68ltr9ljPf2UyTNP5OATpZNz0zpOj9gk3jqBlGGW6X9ks7Nf5GmuFEcqggJf
rXkuVN1HIj2RTv6G13IfelWy0c7zot6eBM9ScsvGMnacNfKVvIOcH8uopH805GJX
fSTW+wJ4COVN8bLKjJKgvt5n6fqTUSSjtMhBPV3dtDnxB2RaRRkaiHIspR8vSYV6
boM5bJUKgqK266FRc4MZt0Tm462CFW1IaSK+DqFgKebWauV6JubPifEp1IM8mgA2
8R/GW9whNMZQESk5E988phPBE2xL5rOxI/DXDbXYeOE5IZSw4ASeGTl2n+QouvaU
EaLe83UBsns3EDDAXxPVxt8g2CbkWbkk4zH+s+WdKudQBeTrZTaVqbK3WenweIHT
4bbhKnjYdk3Ly/zRkdTSnHidKb2/5ZaCe4I52Lj2u8mS8Skg2npMnCJeRxgBvWDw
f+yzR+eN6aVzZcfWlLyDQZceHky+MNR2jwkxYigafINYueR04T7pMcJH497wsuNM
FMn2b1PoG/FHMkQmAy8qCRkkQ1DRWkSfOWDck9F2WTFFLFozJ3qCbG6alz5xO1q9
j2rqD1r03dONdXOMleQ6rfff4EtfCcVLFJKULByA3DehfKrzqvIKTjLKCGv1Z3LX
8riLxTjFOs5V+MHDlmHwiifcmSTo4JgTvIlU+CYJ7qrC96Se5lwcTvfnwYgr6wKM
Vnr4ckuQRxI3cfga66M2OaQOrbx4CiKlO84Np7f770WHUtWC8ybP3t6oskwiCgKI
yJkuKkppTgpPEerSeMMtvhY7OMmEmq5idNezTiWldQSi7idqKqJEkwkUTDut3uS+
+x8x2M8bw9wuijNBnBCRaVKQAMUhj2chh6DqtCFz2msZNH3GoUE99MoheP/51BLo
zSXlO5pEtFwOd5FSThMYE73iAlFf4ic26EMiNJqeq565hkovwS1W4Nfhc9hpYuUQ
KfytIbCLyTvxPUepJGfgDgwMmrP7k44IrbO30LSW4wG89kdqRAt9aUGu0WnX5g62
vIPzc/lu5Jyn8h758VoMMmB6PODMZrVN0y1fwIayGwTUMTrKxv6l4ryUqlPj11KT
L5PofWGyq0PrVlEP5j23rfOBrveT8wH6011TyaHB6Ekv0Yg0Hm0rup7Iz+QJdv0D
xipUsibeDz1VXpmV9C8VJV3nyDS6F22hUe6z0eWt16+Z2lR6vySQSyewlXBlm3va
kmsjLTZg0STSt0JWF1Zu3UgeTdoiJgfnv3NYk5+RnaghLB5EYgUZDFTh9TbAnMwU
G1JQUW4cIpoTTMY+Da+E90SevCFMtHgYwUj/dnp2m/KnTQKgd1bT0pxHJq6uERk5
kuCnkFiEeYi1aTAL1/2UBIX5E3LkeOBEsMQTrLD5xYGzR4W+fSXFvBy1vAI0LviM
8nkbGV1KFuonog/ANNwp2eSwaRzE99CMA5jwdCIGmxOs0XPKukbRGLwa1O11K6iM
QkfAsGSLyt3oOweZQLCeqdnsvbptsQQiWutTWRa7S/29NFXJwBd8erDtmvhz5E3E
qi9v2LZPzW92uWiKm/5xCslAge9g7Bhz1Se42GMPtqH5vnHwmCmHgBK2Ixqu4etG
0sb5142rNRzQi++yEUdI6ddO7yB+bR1MhRXdPWLB2WIsVlFZaQXCTJk25FE1VXQl
MM/ks23wc6BRzE/vrRsZI1lm0DCssOXWq7SW5Tw2dH2qipZiS5GvYFrcHgavzowM
gaV7tRRYrfRouCFqg+6u02NQOZBH1YoEew8fwSfAc2DHEP/DAjWhZnI1OFGAe0+w
GJkIa2Zx9AaD06THfbcYfSOvQRyqkVHRgGu2hAQvYFZH7ORifR/oHNsPBEIN02GR
WGAYe7QEBAL2gTQ1HRczK7GbtY4xgEZzAEVA8PI68VdohsCJ6ikKVu5CfGkqPdpt
dnxjNtcDbbGX265/F0ovZ/KGXwttNHiBQ9gEgFzfzHKm5HjVgU+iL4i3rP007zkt
q3tCDnafR24ncrfiaWvizKVZk3URUyGyNgdY8KooXqB4cvDP3jvw0EHyCIntER91
xFra2RfDobpZHEL3AuMgYCz7kq//HEE3hkbQw3vx1G8sBK6KDvWbrNRkNmg5xIsu
qG88lAKcV1NmgDeZyl5OJ9PGsvmaiapiZlueCGlvSSRD610xzjoD1UlWiSeX67/q
dAPpQzUaWWAMWSbi08KsefK8DgSpMvGG+NyAcgp8fjGnLN/yTcbk+eeEYVAuImfQ
oQkimO7SG5gf6zhYm37n5K+fFJZPO3Vf7ii1fPYvHqFgBfJyxMSMnSs1kK5KzneT
EU0EpzCHznghlTQKrqLUzOVt1+ZVXRP4FitG2h86DT/GOhXb58wFwH99c+w4eGPB
FPq9dhi+FXq9a5fB2VikNubH0wZCw5I79QXtw4WyLi6cFoN4AsA388qHgm8qxNtH
gELW5iQCbp+y4HKrRHySPBXIOFQsA3MekwjfN8uCRwbaElq9vlPPOWTp7rdyi23t
Ab6dCrPez0BX/2JyB6f6YnmIdAGTOOunhTwZPOr6lfUXOXBwQcybViUxACWjJdgU
1rzUVhCNB3SyFcOmrL42fvOLb0TXCIn62aT4XCPDoHkr4ah3FapqPZd+T5UIqP3f
3LbMA1GG/aQ4015NZ5undjC1cdA15Scon3fD3/qqItY16yB6Z3VSBxpz3XsJJlrF
DYmjPBffVUUaatQASfJJavikYpfmrsQoNotrrlp1xjwQPP9Uu2Np+I3am/aTLKNe
k2cGvAjvOuRU4LtoFyTKU+DGVm8QDaRDju15zD3l6FDPysLj2Nktu1TmSJhj3adw
b5RGWDwe2wV86AbFLvMrWKmQWqReyqdghPI+ISdzIooZykhuPh0NjC7NDzxUIr5i
58+Sewaj9KCb3SvUua5ijp8wlZ1JuLJ1HTYV2I9M8W6NWxuy17mAehvcVNv1cHIF
H7iapYQJbcjuf5aDwmgZLfGzEP/JJKhlgjCBFwOYQpmUGCYe2TyvyaDaFY9j/zb8
zWDDgDmOccFn78B67cBlOz2sKhm4RiUoyF2qzOj790LqaRvSugtDrcvd+TG49dfU
8BXTBbmZeUn7soSDceIZLFwzMnDik1xjUWbeFrnZ/RSPguJkMGNHlpFbtHYFEfs0
EkGJs142G9SBDqEwac+BHlcVDrVWXRaG1UIDnntgQV7L/6rOVk/UINpz5j2LM95W
Zq6mtwwLcEhTcmett4XiFmd09vcFS3UNdVEFB+kGwivovRl4ZCr0nCA9VB3teSjO
th0bcXkV3fAEhvC9nJkww455k5D4TnRtp7BvN/ImZ/cqQx606/94o7Nf8G49QPFK
5BhOdEb+UI77s2JqZTh/5WtMOFXILepjExcoj69FZ/W25su3MbK3LsVv8RS4OzJy
Dn2xRlM/gkdKk4Rmmo7f1nN/Aq810R4YYdKH82UKbueUT70UCuBYOdyXqEdXp+EC
f+rlBAQNj5nSyYXt6/akIHrUnYgFhdpJsboD1IkzNewrYKmA5ZofZQtoZWBdxBSx
jvoaAbooPHXuPELcAxzoeR4R8muBwZbe63j5fGCTGz/d6L3hVFUDZapUsJzkWRul
YDzgEW/n8G7X+wixAl5cIPtrpl699FdLyE9aBHqDztJ3YUi4Q3yqhgaS9duyof0k
sqm8Rw5pxuTteg2CBm01HnU7RHITU7Q8Or5LrhceT23AhqnZ5HR13Kn82jLU2/3W
cj3gVKlqmYY5Fyag2VzZgmcTQO++pfOpi6WnVExID/LbF6fd8T9EY8I26ZFV5HSY
3jv71+QLhyhmJxVNOWfFX1q2IU9uJ5wO8SBZ1qE8InBiO7pBZ+Xx3XTvUZxyR3f+
Dt60z5300p8gsa5cOEfAQrDHEyxKVuUkIaciKBVViOyihh+8z7njuButzxMzMwQd
5J6RV/Z3vaZqy/RcpjedWnEqmRpcfm0AH6KLdxEYzk3MeTG+fb3SabT4pAZGx0+L
PCCv8CRT1i9yfks6buGdeufAEfqMV7oJCdilQvNBuRLZj8zvgZ9MMFSrkX9w3NnB
vp8hAHMbTrM9WVNeFbdf+cF49mF6hZqEvrPQSKiuRvQWmM6MviTk3JpH1219qsqU
kkaS4FSWPY01cnZ7bpzuHm+AWtBOjPOLMwP8IOpLlm4yKRyCcHOUpsZHztxNTCzV
kZq2XmykcKnmBNPzvaBW029cFYV2nSt4KHKtfQdYykrqFKXgZVFy196XAmpzaMP1
AtcumdPmyCPsjEumUICx1bWKUCIZjfvgh/oN5DNJ/BaTPMg51mtUCThM8EDcEGBu
BCqEZiyDpj1UkeDtAfu4K59p1FPRzDbnn6iHn9fb4iCqXueJF8ivadQ4Ht1iq9e/
Cb9p4EH9bJstTZ8O9qzZYhtV/pbrdtTXhQBbuQhv1hh9ddbA1hI2G1Tb5ldJdypT
SOlFyy0ttVMSUgjE+1U1Vn7VL931fDgzbhzBF9DbTJybTQ0KJJPqSxz8r8sTZIhl
yc6LLZwTNv2bz+fidxfAhjWUr4/reqZXn+bhVqQgPv2NtSxONZT5ogRbPhlBJNf9
XLtlXr3qxSRmG1H5SfW9fhAfA8UiCmAUJMDkHO3T6bnI2Yho3IgmdFl0hheQxa0x
kSDyu8hE0BEwe6/eVOVcV/rqCivkaw72bkXB9IbL02VHEhAn+SL8VNWmuzuR1v90
r5xb09u9gKb5mbiC61ARdrqdTDqKLHKWid6vpJyZ/KqXTiSu8VsfEhUfKzKGM1rs
7/3dgI1eS8dB090amQqXJDPIGu13PCehS8gSg6mWhX1Ma2Dscz28AbJkgdOn65Xw
eqksFP8CHX0/96z2AJIEPsKpdr4PLOT4Xw5HNZVBjvULPfTdLwPmD3K33yRMLzxX
mm6V8r8YT1xQpkV3Aw4E5mH+9aMN3Z7TzsRYSRzpL6ZJpz1/9lYShgEixGADy5QV
LU1J1/YCqCt1yIPmb93WU0aeY+SzckQyVNq9iue+CR6ZFCmXu3tTYWdcoW/fxrCU
Zc0bZ2EsDZ64t9A7xGoZLbZJGr0rspcp+iuurxpz5kdfJp/dfRBFmgbucn20FwlV
mOgI8IBgUXMN3vwODppu+UZRRJk5P8PB8jGlzH1cno1I/Cf+Eywq8eOj6nAHr/xR
9Irx+qnVEQeZIoZ3f0aWlFruMt2+ObZBvkrk3/QycRnm10+s5o9VyfvXgrFfY+kD
KgT4y75DZTlxWewLZVF9e1HCF6LqupznpkS+Y45Nn6FCdO2/+nI6MtxJNA6BFZWa
czFqGVW2UmwW5TRVEoCbsqzhSUUPCX11mpxZ3M9jHRivgZMy7Gtr8TFRUQ6RShFt
DfhCbdFThV4+8xaFhqwELZlemq33zBekiANWip5fNcS5gtUuy8pZQRlkhN0o6JRs
m7Y4mTG/vxDGClJnVXTRahLmC32nt5JzxKpisX7JcBOlgb5WmlTQ2gRUdK4WMMvt
VHjomDgpw81deljtNzEtF0H1d0S5oh2YSni49DFtxspCMRJeYqEzD/MzKa/1DZlG
5EM/qRqWENSerwslVjmFGUuaBTVFOApld5d5n/u6Jc1ErXeRaEi8JEo+zAxu8z5e
hsatljc6i+BCWxtBEhcB8i8amQYj/w1FSSZ3/jiz8lbY77N+xc9p5ipQalizSvtS
J4Ld1SIgtw2k0MJXQ9YOe0baw/aCt8YIua/Z9uz1cQrfIxKiIXQuglsNwxig12oL
yergoMfPqxL7UYEKOC1dt4nXT2ATbC7az2zxcFWx6mbVRnF8gOasFSzNjRK4n1jg
a8h6BoYaP8gx72r9b/eONfHDEWv42lECp32r2yRm5sTJDClnDk6ZlzHksIsJE/cc
7hJlHVBRLndd/jlSK85dl/FAM8OJyQso49ue7QAIMvmOMpMmMrF5L4wHdWuUzpka
vVGF9dLBbA4DvCga3ecXpE7SPv+Fo10qtXZcLBZWTmPfW1MTXmq/9D2bG2nwOqj/
9++6byOnr9Eqdmm6I68BJGo6/rRxPr2LF8/Qb3Oj4kL1Jk+mkWfmGa7TvfhMLidQ
V8qeCWPf/dD0ldnpxSJEaYWjYd4HWxeHJRIMNV3qh2Te/kllkrGTESpxWADrX8NI
jd8qAfPdXVB07wvKhPJfKGUpKD7UgflqYXhtSzrnUJK4mUsW8Glr5nOl0O/fY+yn
kUNuNfnS5KwQfq9D2dFnsETFmd8JMHh1AO38cOhiFhtTBBnnPqXJpu3TunIIde/S
tvoDKXkuASg8QLt850RHljG3/pRy/e7D5/gaFoVRwBCS5HHfidu2NFrM009CZ6BP
9e5BVgDKEydXNu/BQaRp6TmHW6bsFRXUQape/ALmFavoLReCEtu9RtEbn5VWcxtu
fsx+0RJM4nO4vFUFRvfzZLa58CZZBsQ0G2FDVpqT3KXIfx4eV6xsYTmtlatXDI+U
15cV8Ce5RUUlPgjFjshl+y698yergLbXjqhJ49RCUpMkV+P9l/2MIOWC6+KZa4K9
YKGmfY/Bq1GCad7kYJJF/MlpCxCofyvHZ9AELEDAQcWtJK5taJLocqYDyWvZClog
kcZ03IUJgLVhdLPgrDqz6LFUpQeI7r1JzczMy6Ic5+J+gueDUK00UsCNVbAjp8Jq
4tzS+PDCvmu+qZtqXF8Hum9BUQgZU/WwfGmFRQyjhsx/8xRH3ZsXtD2K0tSEzMl/
lg1Cy32donThySM8jc9dGHVjWRQhB84ujAaLVPhyFlHsqCTRN5BizS/M9EjnbhbZ
0hxqsk8wfKGVAnaHAghy/xn+s/B7JALDrTReOCcEOB9rKNtCm/h9WQepNfVYnhdM
fFtwTHB0lKmWu1dZ5xIacPLtu4f5Hb0eliqRrbqo3X/2ASOVZJBE+zUY9G2PGMaX
JkUvAwyd0DCzsIbeC6pMC9V1asf2wCgZu1KEjmMsdOR+kwAXyzhBCV4phti8WbKi
b9E321TTR4JSIgmApfq0mFGbVP3tLNGyJuLL4RX840ExOTjuP7w7Hvpa+tPMAU4c
L+QZewDmv2bhdypVURn5ZpehIQqYZIAc5Cxa6OPnpmg8DssF9A0lsKgv2JaP16rX
Ljv/A6OYheyAjEdtJMX4sukD/esOALuhOareUMUMID5SuNErvmQz1wPCUBnWTUDl
AFPTWiHu4L/SViUxRwVZXBAjmdDNRxarDZkj18p1P2NDj+py1UJQl20AyF5zQRJa
vrStFmtx6YIwLNthNkukndzsipxQCVKmYxY/fChtuuwHbPBLdYz5PXys/mWd3ZBJ
ofdW1tVeBf2crHPUxELrgVBPFO6ov9hWag5NrC0WA1FyhSvMWJnRUhmx346KPKJn
D7aMgX9RbiozuOn3Ukzlzq/nk4SMyTlki7BRfht6bmEJpzTyHQNwB49PHxqNS/To
M8yyC4aecOJfl/Avx/zL8DeQftEi2if3Ee5K5QHK1KWfETCqkEatHtqLYR6UEJLO
139PPUyW/HKsI6yZqcddN3jSP2+Qr4EbJ7x+SzZy8q7NNCKaKXcpmUc1VoP3XBdz
WuJr838hv9GeoAY1W0Cj9R/7yUjISWxtxVU5QQiMoLVhU5YwUy23I2O8ZQTGN2z4
8dtU8XsBJ9u1V764ZV7nY56fRt4C5tpZYzhAE+CFm5joq2kT2jnVkKchJ0Tgu5Lq
4lcbmu/HBXQGvLzJljW58kHG7qR7pio/BN6SUJNFGOpi02bqVXyELSyEEJoC4r7u
Y6r3WzWu3uZY22luOTj82da+OJimB2J0IHZVixF8bJxP0UHUU+WQhSSFG/4kJJgw
C0MdxQvKyZlm1/t2Tx5mOgZ71tt+R8yCdcUupg66eY8BwHKRg5iPKOzUjsdjE1zM
4258Pm8c1TdLlieRoTynYkK5PPHXRjFkfnUghqATLEllhQ2kLqBEOBJb3MxbgtL7
JzU+RnD4eBLG7khcH5KZsIY8ZzZCkzdi/A3JcqNLlyLLEanW8Vg3B82Gm8OPl5CR
2yOKPp2mzWV1NTU8dHfFWtnAmJosOprgD8n7LnyRCBaEnUdq6OjNXD/dK2NG9eGL
GuV9XKF/7EYMQx67jtScxYpoPbYO5CEcjN8YXVQaK3LplYF7/pVsmuf7wKthpB2R
zc+WWUMidzAUl3paQQo+ZSLO3Wbbzwt9x4Z8sZaVjIwRrHnKQHy6MpKKuOhTL6Y8
xlaEZ0lrVOI8gbcbkSYL0ZiuEbanp9FgyfPMO34TGbKusiEwZLqiZuTZwE8GHmTi
HmDpsXr7DanxYlbp1+lc653sFZnJIZ9JFMVsw0YI5Q3gBQGJ6NS06wki8dAOEL33
bmBlJwTzh4kxcYREHMHjNXOx4MjCHYEODIoGz9DhO1f63KHP5wtr/t/C2bh0TS5s
ucklyHxxwWrPe9fNKcl/FtFKE2Q2bwn7uKnEG1DOhXLdsD93ixXeHwCQFPR73YSK
1eGLk+ChRCzdoxZl6u7p63BGGOXrZkiHovsPn960G4cVP4rbH/gfidoZOvcno0eR
zJWA93t6HJaz0yYwp6hMcJX25gyWHRWr2EhL09IvVxPCz1u2/efQbyxjvBZ8Ylbh
`pragma protect end_protected
