// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:15 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U6eahCnGCfLJUgd8YHb2ylhKpXHXv862M41wIeoD3tPylP/oiSZZ33iryRDsgAtx
DOwCdk0p1rOofy9zhNr4x4vRBGN/k+PRyKREcsQJJvytWxOpi/zFwBD8RhKuASuS
/hP9eoNwQy9jsMrvI9kxAFBUYGpJs9kQw+3I9Yc4RDg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26032)
FNPnr9VeUanqvjVVrrx2+8X516Ycxr4j0XwkbErwVn8uu+MPgFQw4P9WqudIzhhG
Tr/JwtMQmwhOisGLs3b9trzMDp5+4VaeMUxmqA9BgzNMlm19IzWS1qJUw2FeG7Op
UQyWqyVOIQpk18XY+sXwdHqiBLVltwQ2n+vq0BrhwV56L3g7Sy1soTbixffa8dvJ
bJb4QcooeRPtxwM8I+3U35RyjTgB62OhkdgyKmgrwD1lRtfL8fv9yOON0/tzy9AZ
tfNT7eNxkxMTvmCt5wqvOmikc1yOgNSIlR1dq2BjdUqMaQTKDr5SX3ABk0HkNvwH
BUOZBm+YpzCbu0oxSRBk5ZPKL6VmHuf/NmZW4aCCXOqlzO6TC+hRuCh7sGQzDL+t
vKWmrLaFLzLcMLB1skVMCFEiUBPOpXuDZoRawqaaxqTh3KT+88peryY3xH/vVVJ9
lG6uvEV1vJvGcgNU7dFKWocynpQmtqCcSRNjJM5KyF5Eze1kS+5diJCoMjk37vcU
QCTrVItmoUi2SUgcloKrPSMWwu+Nl/w5JeLw+CT139EMMCTcN4TLbskZAtdnDgy0
Eb9RVZ538p0FfUWav6IuGVQ4Z0WirdOJNWm6F+ZzA7bRWUQ8WErDqOP9atywiM9e
Iico6Oryd/NrZbUQpt/WXiQ4h6Lz7SxHCEq/+R5yUrqWUPwvv5wGjHCFC1dj1les
3dnG5rD++SDeNV1yTT3+zenFaKKliLIRwgSW2Flwzb7zaLiNVbq9qWOEQMFFykjT
mFpv1kMNr1jTRuyGtyngRpTmcViLdyUQWQWtMHem8kh/uvDc3OOPbPSf6Kv5mi0I
J6ta0+EhH7u5NmBi5ADeY3y7FkiOAMY9mO+J7sYpme6ksy7KzD15IqcllfKXjxim
0YpqO16ZJjLuapND/yg8WOz95WNv7MLkV9lNIJ7ISiF6JuR/16QX22UbmIDHqAen
AbuyIUq87Kz5WbhlRd4pXtoMZpwIOZDo0aDG+SWsohEF6C6JqSXKXsIFblq21XNT
WyPIC0zn0gc/NW9ZK3YMMnc/e4Yk407qMLG9o16ONxy+n/aZe4zRbgVBmohZonMu
78mJIV9xYQVFMrfO2+ymZC9vIzyIUVrwTOBMOkMxc+T7rYNBEtGeqaWn5B0m+nYq
L+Sk73BkDK3JfOC67XW6zT3acpHiLSGGnPdjEtpy+oxfQRzVJLEp323/SMivCCU2
ZxKIaivCL6xftDHIkC25CXHN9b4S5A7fG3Qw23feyzT0Ji9KVy0yistHp43Je6lT
h0bXWDmsOjYLJP7daFDv/yj3ff7HmlHl8PiWCfmPDN7pqqn9s5A9a7JOvjeVlE4F
ac5/uL/G/Q+gRU8MmJPEuGP5d66gV/mqsGV4Zj8H3Jj1SwAEXbKvUAZeF8SSKHuC
lzhcZYaI11vkNbyTw0FuwmROHrkFPvPP3rdCkvLti1V8JZEAYH/6nvrMCEC7D3xz
YVnX7N17yBXevJU1kccpPyLX5iDmkfEw3DIVZya1o+I1A2kDBUOZT2LlzqGDD0vo
wvPaVX3YjEDuBNz9PZJd97XAE91qDc+8QA5py1PjxKU/718msC4KQT26N1yLKmPh
pas/bJ3xBGkpk+7umvmQJIVCS/0+J6q/Tj/va0eeW+LBeVSQdWLuoy9+qCWGci5g
pjysUDd3sO5FNS42+dsANoODJpeCTIlSFOya31bB8URYcCN7exQEkOTshB4lJfaN
eEktGqJf58s8W8r20pWRacZdRCIrQhQVVMENSkIX4B+mFSUosiU1ZITYB+dnFiDy
F0aLbl+n1BXrVYztt5T8I7WOULmiOGjHN8oSzPSrlZUAtoYNULekvJmG8K0/q9da
E+t0DjdsZZp/l2/wZiARKFMg/gaS5gEYaeU7rf45oEU2NIXam6CooRQ7C/ifCI/Y
CZMT3jgTVE/kCdVaTLneVDh1n6Fob/m7RbC+Xdtj9OYMayEz5zZli6Wbpxwr0P4g
nf7QejiLlvWv0T9EZmfIbvBFAa2wcc2MvGM4Lb3GEeMtuQgBwwdm+oQXRFuAky9x
dP/Acte2mOdjspIoOJY8hnqEyN4gH3bZYGaVK+S40N2YtrWHZvcCavdnvw4ot2Um
/rK00xohOM6UA1FbMpAiULYutPYgh54O0fJMhV9SHOt0fQS00Y1farDDdKsPHRzd
k1fKkUnmQA0g9FwC5peBx0WFmbn1WvV/JmeuTqwU2i8Y8/I00dkxnBMhdH5Lcivz
kwtPLKJPyPZbPrP/9Sx96lREXpkTm6qvxxz57g5SRL7jkl3JTxplXtEvvrFTXS7r
tIKK34+sr/EACq9KLpqAWhZPSX1a7jrdTjPoMs91IFfTZEXCdbD8p0K1UWAaEpOR
Y3vcHTCN122QXvszdI24gymCIG3Y73PE+ZLBZpSr0M29yB8/C+IJVWfiaAuMpDmk
MqOeiTwUTWXzQOIPdwatUvgvYgiQ+iWq/T1Jr5XzBoBP8TyR6gT1Y1I3zNb4r0KG
xHQNyea62qMxPyP3eAhlodE9NWJTzgn7ahXimFQKUeSmehsxY2xPltXivvDrGQ7R
3ORgQNfELOwmDQCvNXb8Y3JmdcSKJNtSIyYgZm3bKlBxHVgzU7zCqrrMoBYKdtBI
qOzJG3ILW4nv3KobvPLfX7AY9V6nM/QlAf5SqAAuNzdhxtLxEUpOPQ3dLIL2wQay
yuXEhoNZGz1eGdRbZ4E8fO6dnwBdhWHI67zJjyeqiuVgixljm0oLYnVuyX0igOc8
U6+u2BgC3iDckueUFcGYuQVBJ+MNERul0aDMhifAgaFH0Jya9lRnjBp+zjt3hVNe
iI/5cELI7H1bhtWbw6nSA9O0C/x4orBGUbd4WenhAkiY8FFygHTmrBAqOCEC+EV0
YA8mD8URsw+ysLe5hdkxHvOPKogws2tHUeUrF6UHel+zkCwhfLk1OXtTQXpLCEFC
F8bUDZUI0m0cgR6abT/FguFDAHt2H0VWRP9889c4jNiAfugqsQz1G0VB1xZfeDA6
xdthb5flT25Id+nDkxui7E+jGuFQVI2dYlS8NTSFB4w0v0GMZGGT3FTCyX7bJD77
kTqj5r6RHhE7uF9buACiQk/kongH9iv8cxxyVmUQ+d1gfxfdlS8Fff0Xn3NOi5eH
1RdcTF0FQoyXed9RdTvTj7ZHfS/Jdwi7U+XxCXiiwR+ruyDfo6rOHNiIGfkrzW0Y
AS4tPLCTsLRQiGOFGHFg+S/JTaaUernVfsTkTd2CxCSq5/bVpxDINLcji+P40b7Z
rXBbWAvle+MipfuPCYCgFbcGtaqesWrfDs3/36EmJ2mw5g/DHSjBhCGHZnO2JklG
/y9CTWunefvcjK2XVVjyOJzq5EsRLuS4CMGJTr7e9tMvjxjFlaWJMEe2/caFaQxe
Qnp1KFiEfVpHJ425QlcVpQNzC2EMxULcWhHllYvGANIBD/GTlvVU77CW4mldr9MI
H3SZ5X679iZP+6rcVuEV+/4qZtscj9l1ltYHH8uWaIij/aYaHPaep1WOCBZOzr/F
rmWXIInySNskaxCAoTLXv/UHoYr9V40DlVI7KxpkRpDESqiqsUoBlBPsbwz11j0i
wz3SUMigR1ugtCqhMbII499MDYz8QuxHsKYHK8jPjO5U6rMaZQfQm9eDWfmEGzeK
SL1AX8hUeByjZZTUlMLk7wCMs4nC2kei4GGcl52WN5v7qOcBWVRdLmvC4jV4vn8Y
dowTDt3BuxtMdyXW/FQKdH3vqpWqRJZsj02ojfTamjH2G+D9ENcvjhC638/vQ5zQ
7YauKKZD/mzQebmpiUzbhVcyMg/dwFSDTLYjAYejCc4ekXdXQrKVjwHiWl7Jh8yU
DOfCuKsBLU6y3CktOG9JI7DEhMO0kXWwH4dJ2tTWpgk8J80vmTZ5RcWbNZb+nKs7
vYKl6VFLRNfg4R0NzWj+zij/wujYoQrBZqKvruVgjlN3+NrhA8UVIshE2Eu0067T
UXQu70Ube3hO+ddsJ7vb+6WAXfcPTJ1jdH8ge6OFTgY3rSzzfBRqivl9RuPFsAnk
xlLaaqQsNKFeGcypXBP4jpfLyUXnl0HRl/7zrFwNkJS4+k8bAYfxBbre/wx/RA5Q
dHtf5n+MTLCgP+GTSSWchHjV1s7N/zj/f5k8qDZIWp7McJ6b2wfFvpGNBocdfIny
c7AeoBAFezpuzFF7KqbQeCE1yk1S2KLeJ8ZBWS0hQjjWEKmZGNpHPOnb2Bwxoz2i
H5N1+x4A+bvTOr+pRMJcdP7h9ecVEDKY8IloWFmLTj33G/WslUfgZ3pl/esci1kS
2CDYrzpQ54tyNcGq4uRkFqE94PxFEO/4FrYoZhvD98uRmZywCHovlljVgqYvKDiP
hlViz3SMRQpvT6Pngcnnfu49V9ae6Bx9zqKJ0CZHFStSVNqazvmVaDcgsx69p4jc
uSnP6D4DSpvX+lxYoN6IKiMoWSVkREQqx1EBE+t9Gak00xJDL2FB1g9P3qHOeGxa
mrLslM9aDpmMiP60TpV8zZxdcJAKE/ZR1XCqkbKt8SnpBX7NXk5Tw5tvBNUO/tU5
yukbg0ZI4J76WFD87Q6GFDOnWlE8xCCKiSkTlw2NOWUqbjfBClbJH+s4YK3qArwx
y1Hpa1EDsMTMuqq6Z+40md4gFd0GPSENNSoopFJR6aBL+OgtseNc58qBpp6QK8s2
kl8LHJmkES7e63dPXh/vlhAUx3OVq+pQRpJItGWzQWgwgRFlevPVH6SRcTagU4Bx
tzoEpbtg3LFLFKgernzeNfOLgBIze3EKzPlsNLnZbRD2Dd6ZP2lOWfdgNEyo2qDT
5Sx8TPR+enXr44ZKGOQEfTH/AGd2ob6bElAW4GVApf4+guZ7uzuFeJC9Q22PvN/T
KyZ5x2AAHuZ8ufWXyJGasijcq3r+x/74hhSA7oQjydxZlJMQF71mF0Yw6vW4nVWj
bULBhhHy5G3rGedKi1KxGeFEFok2/CVvcd115pq7LW40ez7QN4SwbNPGlfN4lzGc
DsVyizNpRSrk3QDVGMKVS6FuLy+KFSaeGjGqOgyqdsHEulFEqb3mBUYDXMvlsa5d
ebiQpTp0txQcBdfK0/6986Eli+QZPwy78XUWzXnGmAApRaMMRhSRXJlR9DY/sui3
h/B2TnABYsGZPIZvEoYC2eHWq4eUeUfQbw2J6ObQktdq7tRrbAXPjG64DwAQ2TQ6
1OBlpp7lJ6P3lrTHbh413cJ8avBbMG71b8VVusS217mrB945eFtxJEaXhsVcW+LB
Uzxd7FYYJ37DEs5gWRNt5jCYBL142HMpIEG+raYGp6LfeZ1MvaxYyArbcMUcHQG2
PeyUAPjk12GR8KandFoBpebaNoHMRrKZSwNHGYr2e1D8ek16U0BJJnKcO/Bqk6q2
RVyYn/DXWPBPxHv3PiLoQHLU20653uBBmvy6eIP0/k7TNz+fhOzbMA57eu4lnZ6k
+EgtRpbjdOaFJjwRi7tLuUxiTpyBL9Ibojxhs0OJFj7x8eiFNZiLF2USUZLBJMf7
ULiOBWAXA2AMFz+UEcXKaO1dC8s367XoZPxhyLT8tWECmv4+26pPDJyS7zxZyK42
wF/H2/OSN+GvL9yZ3ofVtp5OYT/sMcwacp2eOALnpSWDZFR2YDdwsDk2ClTtZi1a
IwcqtgnZvOmcxXsRn54ckygj8p8eBlvzvqB+JN1DFUnGBkHMgtP5ysGEh4jq+3wy
6js/HIRUwZ5qv0j3Mz6u3gFdyresrmFf6m+OOp2C7xwuEa4tv9VOEWTM/jnBH7Ps
brkjwnJ3LG1/pfXNSLF7nQ9O193D1FDVSHMFs4iO1THb+8f1Hy2I3LpQih14P3iG
YtGFeK0OTl+LB7qtdNZ/ptxXeWPxFMkrb2DVhdb9t/ig3Y89Wi8PG9PPUvOb242P
ReThBGTUIaZZuymvienptlQaJcxQaE6nGxlJy++xyNwDp8DCmB2l0/wUtRF3ZE/F
2AFwm+qgyXPDlaj8S0Q0gi6XbnhtK55ZNTOcyvIGTyetKc3U2TIgCutaP6alaumL
w2Tx8iEnK29mkTuds8WXcjQBdxrRusY42Sc9F785hSUWrw2yu63kK0fMS0Ka92Rg
zNRxC9zgzjKAphQCnUiNibZ/5iHyDfySNbn4GoA5r3IQO/IRUo3w3p2bbVbaQymx
I25jTMtin7qthQYizLAKaY8XjKhhmoHC3cQK7L3bI61xS5+GZzzVAfnYUW3vhOox
PO+jDGu7ku38SLN7WU1CtbCrmIyMeAXFHxNnwxJ5czbOX3tBlayq/6LSoU2r3jGq
z8iBrnRJ4CZ1dI5XQus/k/p6i8U5d+3/TmF+5Iw2s/LUACI+IF1ZK+j69N1y39OG
k2mXLRguupVIqeCKey/zruJ2WiSxOYyvEdChHD6HereUw+E8LQ3T2POdfeMjWFJG
fTighqgLylv2jHKr3gUbhpVYGbNILw0etKj6u3Q8EgA7CaTntYpuzGbpJMy6e6Ms
b9PbJKSmYGk+vmh0/rGVwFcRX8wSseFES7++JvkD4o2/iBPO4AUhDTSUSHevOO+t
QIcyYfd2BgPEqaCs5CW6cJHRBuTsn0Mr/PIQhjYJpIDVqc73Z/+wLkRSlY15ZTHW
pGXxejyX4MjBOvFkPPAvNKPxTmJ0dev+bGl+zoOJhOYI+vlm5cLLEn7J24wLXqGG
Plgw1NzjR1hkH9NaO+fZVGteD/t2RhXYcHlcRHZGd3zHfENNW162Uk3wSAk3aV8a
8lfhRfbWLlqRCJp4JlW3sSY/iWlTqr+HTihHFmUuX48VAYDfQ8ldKbKPwSQDKZhc
ZzLJScy1AnhI1W3gyxd1OQPA5LVQBMyf1BrY8btnhNffvuTqurCnZ/QdaPLbCW8V
4Z5LwD+m7Z3PkQkU5/3Mgi+f2ixzSUbqQ0UlSTrgQkFKrLQByR33BqEZm4a0xfj/
w/M0k20xnZX4ALg0JDrYRywhuuv4mIp5UqJY91ULnP1N9loKUYjFKZq76jyNzCXK
P961gywZtdZUYg2lx/tmydvCP/MBQPu2TIAhgjzFUB9r2M7S8a/GuZgTmJh+nkaL
Xkx5/6SdmIXRNxCHfW3/1gDUvpgfL2bc/O3EBCkUGhXi9DKt0uCYibWOr9k4LmK/
8a5+UgSFTgNb4MdOQETpzjyR/Sf4WIlaPISI6GZRnY1hZd/xahHqRXwUvu1Tk2PI
8g1VJYs1hF9Olnh1ZQpQLtVb+71zbjJ+BqMpkdeyd+cptm9DnljeU35JneuhDG+y
8NWPceQglDF3y0/I7aRYsqRV92hqO47g3J42WV9sWIQwkH8QfrpmogRhhf5uQEGj
NgLwbWizgpG98kl1k+Ci6sETCBg1WdNXEkmDkGD0lWKc05khvwBTWVvF0ffZl6pS
ErdpsgSSCjXs8M48KHoYNJ7M+hnUVVmCLQVmuV5fUwhz5jtiaI6nTJ+tuK2FGvP4
wGOGA1u+ejRdfK9pIwV9dUQaKal1+2VEXRM60uUmYKijVK7jgnEYVzd08Lezbvno
Y+N0owoUuz5f5rzy+nYxBuNWbQZbbfls2eZZYoW9jhqCsUXBKE1fUafV0Tu+MNP1
lhhrcnBPhLuz2kOOwo9kG+vmiIdWibiumpOy5NMzcC0y9CUjT3cLeslS7l+/lgHQ
JHI/ufjdApZior4iALkDdVsllaceEGwkHpl5NRXaqvasUWPmXLpf5rUDYNfMN77I
MzOzbb2LFRqYCQpqA5Wpf1Kp+L2iF3UH7CFiMXFWowBjzeRZmBQrDT9iR6F9Poam
vWHTuCk18zk5VS4HZ3e+P+/osXmgsGvYHxV0viC8wW9506+WvQkpyuoo+cZNJp54
fEqXd08/x4HI5cQkD1fAT8PbHraywhqNz4waH3sFIMSzsCLEfFohcfjxZdVX8JiC
bNtZ3bRkQd2+ohex0MgdVdXjUnpn3ikH6YgL3hvXQDzvNTPbDrTruolzsvJByO7+
KV7PsgNNr89WUEdIPfiyNQ3AhjYDagAX4StK/40ZfjkTMovZOKauHsdaVXFSdzKd
yzL/ppEyZ9zIACSUNbuopqU/pguE2mtRWzhn6q4XxJh+fr35ISAsujG5jWpdvKOM
n5ixw5f7IMjisHBDIMJxxvz3vR/ORDVZIISkld7MRkT3STP34u6ubUUwWj3mVPDK
CNiwB2lF1+hpgVseO89fiBPNs03o0raMBQLyaYUceowtmYuZ5Q48ET9vQd4z3yhV
LgFRr00BqriA0O7VUa8ZuwBG3I3jN4qNi3ZVAN51CaauLCQHgdsy/oSquUNRkTZI
3aL5mgSOjdPoWvhnJ49IoQa4qjmjGhPa0SSTnF3yg8MYtNWzeVpcTYub8nHDY5j0
XGzbeI1/abMwIUjGeh/1z+PF+T1kyP0/dbAOSkOTMOmQJygFTRPJLKGwSrePmYSS
J0bOUz6EAOQHIVxcE139WZg7jwp99EHwp8IHS84748/cC6/VQaR9akfpTcwm01jw
VK9oSlgpPRnzUIpHcZigyFtT96fs2p44v5AG0w9YBnOA8NcPiPIlf9HRZD/KFAj6
ONoKBSN3fZRWa1vqOuVTngY/1I2vpHKK2oUlvCjoiNXJ+JqL2vCvZyFX9zrT6/46
/857iYpxUY4zG16YV5HGJGg/s90MmlrfU1DkXXjaODQQJTe+lPZs+YQLyWHMjzGF
ZDBZFVeb5ZCuv5Y9Il296u1Hqk92cPB8Dr2YCA3dn3PRmukpfnus1LhvnPoldEwF
aEMPuu8fAmWJiTXEgZcxGsZLZjp/VogDFWVpu/JU2Wsxnyt67JCi10q6vrzeYj6o
KKpmKDzzRsQP8xN2Hw6IoM5xe6f2w3PHS01UPmPlDK6TiwDetw6bKYwsmyawxHyi
aMhVKz4gHfmQzFOHiZ2onVPU3+9JUdwkAlQQaLBpPRz/qDTxNSfLqzlCT8em8yH0
CBELR/0WNgtUEMkyZzOgJuOSU5rn9b9M4sdTSS+y0zz//ll+ZpCKvg7OhrW7t+o7
7cpZK+ZDw6LQag/9MHvjk36HlULfA494MAuHnXW7Tj9sg1eQ5uHUigZYP8QPbRMJ
EtKHAwvP3PcZDY8o4Pc9auDN33rhXc8UP7HPCry6ZjpoYjBKbVsTbFuPnfmOiXOZ
mz+RN7pSgrNonrJC7qBLUyXJjZw3DHqVdi180AnzL5hRWPQY4H1Hh4qjTtWzPRUA
Di43EpYrykMPLR5+nbRUqLJWwroitBmgsEJwG5a2ijp0hNahzwhcZ6OWFq1+ktuM
t01cA6CvuwlBdjPPUQYg2ivTaymxGXw9WqrA5lDPXa6xNkw/uApkLA0gAqx7d7vR
6/Tw5pVodDnP5J62DE4xWWyEDkqLTfagwzGOvfKlb/Htivc7GHnVvnnYDcoSfv1L
YWPqaxMztxXl33LbPDee3uXpezsWjxAQm5x2hGmIGkakE+6YyLQO2lNqz267DKHI
Zk91A0I2FXk3cqcWh2ixeSM9N/eycfgkigY3aUeCepJBn4MYlb4nhChYujlP/Qfn
CrnkWRgoxiNv1JxgHlXN3KRgYSJqIIfJSEubn+WTh87EVaWMPRWeeZhWg4B8eUrA
RpcSpcXvbKCACI+XHRbFlvS/WJrgKKEsA3HXlNwynz6pMXqYAZknWqLbIktO1qGc
A23pslQjyUhMmLds3rUcoyti7fcwCLfN8qJT5nq8nkI4Ghusr0RLj2rgEU8L3Lku
JEAqHE3dGwuibiqgqqCfNq163MllwmrlwXMKDjfwG86/mT/cmLcmj9WU4VUT4T87
XPCiYHIR6iENXPlOeMOAyC33z2ppIyspT2NZS/UOecjfqYYxypZYAnUagtNphElA
uw8UW4wH2jgCBgA43zNbaStRoLvdMs63ik06flM1096togMTzJw7wMQgV1STE237
YO9TePMbQOgV46nHSTy8jlwMUeVIemyN0aDE2aLVZXXWh8Ah1JMfBKf8cB97hMUl
ca0jsQvWlUk5nprjFF5IOxC+eHKQQWD4YF9sKHMx9TVDrI6ST7E6zmF5fkxuIag4
I11k45/eQ141P4N/JKQUP7AXdZypHvj7zhd3OBVhqMe7IdPNs/4HWZi77cfdGYUl
M9pUbtZx2ZdBnun2p2QjAW8VFiVIFzexbakm0nsK1dm1nQktUA65vaVcK1P280QB
CUhILHSznAD6hmddufsVHPj1EigDNxQvOUd1LE5sfQ3LjJC1V21tqlMJm1ERS7/x
qbHoUvTHV5NENwV3f6x4GoVLeAylOCwS4t2J01sWRaE2SYK70i1Iv5ePoiWl8PhO
OmreZ/Hso7h4yKohNDm5M2xBkc2GL6eZuUICp/roKfgRjcU5qN6Mo++6mqQBxZNt
1zNIwk7Qt+DBcApFsycowTEUI/VZUSQdJ8ucwxgTQWXiEABcdY55It19UMX17te0
kETdT3FSJ1f03MXiqYqadZ/kLJCiLmwC+4rhRqwNyENaLgz/OqsHsvY4UPLdS8Wi
uKOr7P/iKgUBQ5BFJXDW+/EAxz7b36ZVvj6trt/zUVAzKI73k0T1/QyXsQBRTQ65
q3VierJhb1oTIhj9CRVczp6IKF7k+KZ9JIHbLhFYHm1BySQUfTaQo+SXIvFeJymZ
Yb09L/wdaP582xgPGbnP+CBk8wcVqFYr43qFtBh22VgdiPpNsSo+hpd7S7N5Eo/r
DDMqEgIiu4fzXr3Jq2vI/zDk4W5lUhTvDOMKKY9pe9bEDRgqnvxHXV+66Ly0tSOY
8Yd18vsZZkuNwFPKziKqrVagPzE0SzGEbykMYF2Phi7uxhjC4NKGnDRSJsb6ZVPN
frVsmFDHq4dGArwD1SaVT0Ex5zahlp9/SA8uKmV9l66oJHjb6TiDwmkQM1UbYxYB
n8l6SjgXe2A1fLuDlZ7/9Aa6ZwcGbZlje29ax1ODcsfqY1UMwaKYJtNIbPF+jcIf
7cZdRtOCqbRci2TMvvtYMRW1SDX9o17Pn0w269p9NswuUJLvcnG91AATsHF2pg77
Q/Ix1Nd7hgEl6HnbjKsXW7ucjO/0RS465nBJKjZ6l2UsVXA9/yPoUcuqsYo1bdRb
lXCKuG0n3pYzFm1Lp7Yal0EgR5fth1dOFQw4Kw2UgWyeJqQZYqjGoeTYamnJAccS
URCviZqGlkYvsXMi/UmlJ92na8YSp/852wKPsSb4lxJNqw6BEibSaY9zPSEn1BUc
eNgCMlOHW6cb6S61RSgluvTMBLzEG+Iz4dK9dFx6cT+xRPMIHZdR9TLxoFvjcIt0
yZqh/RYvkc8HkwaYDpenl6B1FeCt+CqKs+kzmB88y0+sIimf6C9AHH83lrq+IDht
CldlTveFdOTDfB6IJel3Aq8N7r3aJUOFt/Zb/6x/LE81H1KrS69l8407EZa4fsrU
spmxdT0pPwGKjasTHEis5Nx0+0m9cVWvg42ILa2dCWjEbTOJ6XXF7YSDxGMdZyQt
tJT1M97hWi/J4U0wyxY0bfENKbreQDr8pTTYExaFDPPv4lJIf/rmXD7NnDH3ZCF1
z9ry8LorsTpLYoNy6vyb2/EOHw+Aw0ekWOxRR1JIKr5dZMbR+KjqbVn/M16F3//H
z6OX84krXbbhTQ9zlWkmMOpxrTlg64Yh6UWghBvUNQEyJpBGJ6owlTgZLlt01gYX
9+wVZpPYaW45tr1wIJ3MwbPnS1s3S0E4u7XKaEozEx/mkNIu6i8Emw94aIbq2X66
xYtKeeVI44bvrQkPHP8ae7Zlaq7qBVkdSc/PtXknPF51zF9TOC3DPyeXPMJJ6HUa
5/lTeCZgRDnUY2cj3iv7eOR53TrhnFUXT2AX7PDNqtJJewOd+Lf3tPXHTfPOmlxo
JZYR4SdqhPH+Tgy9+Q6JXinKFwzPmGivEOB4N03j8a+JPI4SoFNBvCgQMWnaX4hG
IKbmSSNQfG7afsSlia8eOn649ON11NNUJPWoSEB+4GDkatNBvVCj/1ORIgRdIele
RpNvEpRGkuDe7p6HXfj/XyA7ndsbslN4Glh9l/jHrQ6E14IGScnjxjf/nS86JlL4
EoRp62YG0TOk0sFxpTbMxhwJ2U9EJV1ywV3kE7hBltw3O7aYYMjRZrUFulnmUd83
6rx/j8MrCwy7+bMpOXhleQb8T11qj1odCW3EKE3D4OWwyEv2V5ZSzJhAYFC5HQop
53zb9jnPUDeVSoHVL+hbrx939w6tN5raLZ5S0ZfrkVpOu6HrIXesAVmHPblRHYir
oZvoPJ7BnPteDWnYgEPdoMWkAJxJx1CXIjlNhjF/vIbATesRRTJKGQROXBHzHWln
lme84J9sNlWL9ty9d+XwtvyyKL/8fj3gWST81vknUVpBAs134gnh//Qz+QihE8Oa
gBcIbT9DJl0EHH/MCXFoxQpPnBK5Mx1MXePJBOTZdw/4+6t0HmdSuTCbhOfxiGcq
XQBwded3E6hqs2VzXG6mxeiHJChtNYSUTSx7U4y3OjATQpaksi/4r+S7aW/2P91R
zgPAo9JSv59BzA37FoeYt3szYENBlPB1uLhwrtp+SPmhaGRBUIE0lgB4llx4blLj
BDjVjV5Umg0rKgJLAVX7v6N1Exb4huVWiBjjdROm6AmSW/3F/dj+5SCag5/s97B5
U4vhZloVPpoDnz73hQlnCKjV163e/Dw+1kMnOKZambt8lTwqD/bcZZfFC7JP5j/l
AQJ2qPkrwHygB2DNYyYgxRVyhBqFmPrWS6UsyEW9GbrckFmORB7HJdhKQURhJtga
Ex3tEnDkY8FHae+Lu5ohR0EgQsK/emepRHkBrtRkJP1Rj3wYUlLWDrt6IDCO68Hd
x56x2rRGZH+dqwYq3ze1/bMtL2W54AvPBNTs8zo0328/m7V6/yM/oRkmtwJWRd0Z
97h7lJR8I32bj/No2ny/V5rL3LI+ra/xkM0k5M3zN5XXM1Wf8QbmqTOy6ogo+l2c
UKHitRqvssy01zclTYsbdLUWHCmF7/eYt9zXcFjZdPavPvBxVwyfA/wC1Boj5x2M
ul+MMNFku90FXkXGZytm07Bvi43hr/xLtV14Tw6YV6nxow4ijOkAooMl3J1wVGVg
maVeWdwTQrZQdYE64/QhfCnrj2cGIZPUSgq6REIfFyk1JkwdqtIkpkqxaaBpXeIf
jwQ2DjL10Ot0Kq6J3AgOZdMUl4ZVRltGpfbNLDSwShZA5j9fYeeOwQn8oMqQE2o8
iEvTY7KvumZoktUln8qZe//UcLYZVhEO9wWQkKJHrfwFkC9mIR3t+GrPuGKZNXTb
rJpJL8CYlb7/U0wiXAl2E3hG5vo5q+nNAhQXQOGWIFxzFsHUmQPwbB/gx3Hf3z5g
4v0ShD6Iw6/8jaH2J/7TrHaLMpb00jXMc+d8fWTOkThIbdZe6dLIbMNIyaWecuNO
HaZ167+VD0nwsJS9BebnHgdfRWEG1wS80rWgVeOa51pFiPwjXadAW1edElMSQVoo
sWTnl+J0JigC8TvqCcg4Mm30x1yc2UoxtPJfR6eC1kenV9JjMSf3pP8qF4NOvn/P
uuRsapBvxDk56KkewdAkXqoL79mxUSCZA9WExwDaVNR0NKRW7+uX892o8VkkTEKo
oZCe702KmVQrpU6t1nkK/aO3gKdpsrV4ovgg90J8gMWZ9RKO5XeDi46r/etvft64
QKfqKp8xSwu10gbBysenIelAw0GcSHGglJ78ry7VYKNT8UY1YPP/ar7IJf3sCgKd
AGX7Ok+6eT7PxLznMZpxDz9Cb1biuCDdjX6jlNKPY82hHQ8Fe68DccePT6l6iq92
vjFZa1ajkP3bQp9Qhe72pQgu8OM8VNkON93u1M6a4MDBEYmzXuvdVg87kdCIvaWw
QVtl3iB+BNNg5zZke504NqyCOZnEJWK6HjO2/53Rz7U0FvU8cMHZ5lLrtfs3l5An
96DRtGZM45BJ/YvP5I6+6XtnkuX3oNqbBiNIU3YCuyv743Yw0eXfHNhfg2GNnY5g
xXtFZW4XBfulcDouRPaK1C6hfQdUzh8kvV9DmABAtU5qIBaoCwfCb/1O8brvqmbL
hGgX7nkzvoKeh3AVKW741z7svy6EiYB5s2r0nUrrzRQpLoi9uoEsSEr6bETVf+yf
ILjI+0Xhlp0kqCsVRcChX+ds/LBibcKIw0JYdGozO2eIQh10NZx8BfJkK4agB8t1
quIOUwoKDPiriIgzVEvMl3oWc+5ne50WPueXXKmKjmawdc6yM4QVU4bsVNeTGP4d
BFz2eIUbOMqiMJYc05u6nNL/BBqziEPjR4C3XKbkQH0ZvpHuc9awHYuZE22BXWKS
6DY+YYL2b7dZNJYisI4QU8Bs1sO0zbtYDuxik94jL+9vjhwXqtS0ZS458pzDAXSV
qfEvfVINanFSaOhoiBgoYMKd7iOrhss0Igh2QUF1JfoHELk8ltgrXCoqX5DaaESb
hQGq38jb2NScIiPsaDloTKIWobn0ZfRfQ1gn7DCmL9hvLeUO9VmXVUKWB7MsXw4w
LrdfdEPTqPkXPmuSOMvu9p+Y0QxxpaZwXOKXLy6vZhfbUglC/LsR124GgfsSfMKF
wG2P64uhUa+Ny0ATPDnOrqPdZpQzJZr66/ykWAhulxSOqMqo+RoX8E3em6fsG9lu
n/5eLCyZnU4v1BVXWU+Wxbm66XpjiDMEXH00CnZvJxiX6t0K9M3HF80acPU5tYx0
6F+FVS0ILu4LeKPpxG1udor3SwOmk+q2gOhuvoEOY1H6a/gvtHLuyEslOsQGAqow
izmthWpRE/iqkTOUFTbGlyaRq1MBaTLtHCFFnBJx1JXozR5OZZEYi2gB7Ncmy7RI
Z81tnuNPcr3DJiSwJ22KTo00Z0QmuDN7HRjkLseckBXtlq3CXU9eGPUEoJg1Gd2E
YyAhryZvdHzvxD2DEyqChZTYsYfHs3Y1n6KCQPaatUzKrsrRn2ps6rrYWFlANu+W
oEr7zxO7eidua3fbHofrk/rd1Df8LbXtypizDnonkSEGjCzI1EwIP3Ml28/NuEI9
UCbXTI/1z+43405Xmig8ZNnIXm4M619RT3auZ7saJhebkDY2mFKuV1K9PkvKLS9m
EHP+sCSwVIWgtEcpwwIm+A6D1S0X1zA+L8RdFtvpIxDavdS5OKMGFsrQ4PNTAyc/
wddLw2toF7XF1cMOepupWwvJfqqGLETnq3K7Y7eDyNAQ9oPTduUHcPQroRwpWSFK
JPEEO9V12DGNrbhxwslUslJ/Ncxu0iOg6nLRVx34Iqc5f9zYSm6xT8Qfrj9G7p6O
k/5f1LKEmBl3vuyjNjMO3ElmrksFqBje/bMEkW25T4T5yyjJoXAF0/F58SnikhUK
2l7KwDwLh4ljKWKMm8cQB/maQQT/vK6LBsHVntLKCGtKV403iIuhPVS6wUNCPQ8H
2wBX78Qfu3f0TuRlOfoIagHoOBjd8fAu+TwukEJ70nHHBEAGO4gRHUmkQ4WlQUq/
ztUMfc8/60EGnRKhVTmERbVtC0e5YTOVE9laC/q4wSQoEzCn70eY6JcYw4BxERps
q8bh+sq7c9Yajrx5m4fWqBnuIqWxYBUzFxywtltfnDaXPzDnkRCeq3z7w3fiH7ar
EbGiTqIkHvkIdxm7pGl3xJRE72VPDKTsGK9tE/D0Po9Ix5l57+EOYyJ6Z/illd37
Cqo8Nkre4nkOFujf2yz42QKFgZo7N6CqAYqIOytXY7+fvh2e0bJNLjCHKf+CBW4S
aalouBhJpp2B7LI10WON4tg8m5sHfGBS8d8WU9IgpTSH+RuZKPsv4JQaxdvv14Gb
9gh/GEWkqIQCZ05K0I9q2hzkHik/KO5WdZhOxWB8nCFw3C/ltR0GxXgXYkvokUi1
2SdDvPkZnsi0a+JIjOtYwIl49HSXSTeJka5XRG7MtHTLmKtFAEtvI18st4oNDE39
G9fn8/EOBLxK/ekP27M1mbf4uOJerReWSWAThKgPpr5SWo7uWGcfxN8ArZbIFbUU
qc/pFd+GGFS67J7eWjpSguksJZ/Le/0O2XlpYRC5d9wtlDfJFENavM/IDoRHIwj5
72mD9y66XmcqziMLt5REAcRsl+AZHFvibyyBkn8BAL8AK+jn0NquWxTop4tuP1Wm
kK6gLa5G6DZFYiAW4yZayPdEOlw/b044rTSi021o/fMJGABtey1XUurNasThC7qm
+q6W5BND/2rSanwIIHmPV7Bnl7lppRlM7VFdmJiEShS72OV2yOAmwO7gCUvUhq1r
3IuG/tz076v2OmE96fAryEAc/5hxDKjlXso/JhgcKYWPRJ1Jl6xJeexyTQw3rwWL
zWRIkb3rmw4jKrzxF7kaNxmvQCe83mhnvF0sNnVXvsGojY7iNX4tqk/cqZQxXG3W
Uimo56pEf96LfO3ou8l1MFWg36HJ17fpvysDPDYaeW7PZ3X9uzetU5KQnU89nvvc
UtNkiD3845CCTE0EvNhR650cLOtUfu/7zL/lBIxXiob3cmrig5tygLoJfdEcMpPz
2LwVMmDDTY32cv9BmGfEYlyYro5MIXcf8JLj5TTdgYXCONlrcczXWRv99untTsBs
R09cz8xbuPrKmxDnH126CrzhKUNiyr0kzt6vdBFu+5o81TRkW5sgrL+yOfbVBFDY
Y3c5CeNMWKMGLEAgQZH29OOpRLRgB8WTQLdKxwQRHlMnx/27Ob4FTRTXqbRh1XxL
AJs7Bx0I9OlLgSKWaFvegAJfUs7Tfyh10qQdOH1DR+BYuMZ0qPRe7HzxobYW3vOh
kWbfZFSBtsosVAvE2eqN6OB3QGsFDOg8xFaQ/4ozpajilfU3JyIrUUxx4Yo+5SOd
xaHjQJI3AB3y1q11u1pmqDJ8J8ziniB2KBeOvG0iPeVTbFF61BjdOhfqmv22oEqt
5i3fjtXpeOvddRgcfwgFMkkBgtOYIvouZS3wEqsZWaGa4W8mEaq71q7ATkuUPl+Y
/jRJo/l3Y9f1GsN4Rz9n9vuDZ5MJ3NR5ltKiBiAm/FlalvkVST75hMrrx/yAANCZ
8UPZXaSZbmyxFmyzEeczK6dUGpHLJe87Mh90SkQc2+vq5ilS5NXB1Lp/5nBT5+Ia
T3VcTZsxw3fRweZP0pm7YfYsHewQTtK01jVfWvk9U0PaSjUPtdItmgRUBxELUn9k
v38VxD/T5Cn7lDJwivwaBC31zk/iHfNWiE+4wUBVRNev5FpA+NLaO3I0SLSmRn6j
+vtY+JLsTE6SF8QsQjRC/TzxbVH0i0S3CQVSoM9OceM6EcFYS5wmy+lgn/ryg4VW
LR1TN3r4aYzg4tyDEemGyqXEwENk2k102KE2PBXKjVDJbXnTT00o9rCjt7JWG2hW
bH5Iyg2PRSAEyEuQFxK1HypuZy9mnzajz+o9gjumHAguFB+umUY/3E40wn3s5uGG
GHJug1T+wtOGjWSSsrP2tmog7yqqkGMbL/Ib37FOuNdf36BW2pZn91BwVvNGI9Xi
QHLsFDb/tW3fGFLS5aE2pbFA0lolxv14ZDFtmeLL0vX9PCgUvXa69E40Lbqm3ZlD
yWJmrbBpMQ/6uzjeIRW7WFUCuJgyC3E+XGvc+wMIhXAxoPy/JiY7gDiyLU4jQzdK
vu21SRZ0kYByHdHGQY6hrOxa08L3f+Y8tZwwNz6Cw7JBrpQ1+5ADMGrNDMtKTsyX
wLNPznOCIg4+xO0iMKAfL1/3wp9j2py7c2OpfBYq3sKJs6T/NF9JDOjUoaG2l/bs
vzA56nK/hDZZ7Cc9fj7pzYXhf3ENaGNu889QCokibdPi4NVwsXzYQ2IDR1/Dg3FU
nfGwk72rqvJxu2JzrOyvx9vwsDUdm4h2Z0cPmZBCoHbTVEiDNCRb/AVwtQI8xXXg
bVaEKAlwkO5C3nBRt99wannq3MJ8fXdVbWW27z2FVTWlVT2h7Lna0Z8A2yTYRfZK
4hb+1LHHnbKQq4YSj/A2Whggnhd2JZrvBmZaiAPpkDCBw00Vw/CUbWOB3+up4lHp
4PVeMSU9H9HznjNdK6GyQNhXK3f7Mi90unoObdU9fmj01/pTeNgnsaQOIuHEQwBr
5wGqRnIm7BwmAWVGqV/2z5rKbC+WVt8dSe30dcqedRx5U8YU3E1GrEyZz3nJ94Ks
ml+XAGLcmXuO1i+1OdspO2/lpjItpmJ4IGDvrUDjPkqWuaNJLVX8WrFjrlYKeEeA
Nq9XFkCvzaERam7os2XdevDNhoFzeM4MKbjJdcOOhBECrmC7Ewu7T8Z4z7mLTtiO
dtKfHAB8BCq9gqKM7j8PO4MsL6cygTtNNkB6mt2gRIozoJhfWk8LABfVvl1F2t/e
+vJmJfSd6A5llOlBfWudWWdta7R2IQVgNKYVpCfAgDJyURhoxImtXg2zMJ4pJpNI
S/dfw9J2XXBJa4/rnpnx4q25agp4hFflu43coiurNohx7mU+IefT7KOzJyJT0Oyt
VEnz0pMRQtpZIibtd6mLGgP9f7TlMD81W85wPSGjjjz7yyocXzyv2+vnby6hod63
k9aZ2vlqdKlbm/kO3AtGVPVQqUvz8g08d6QoMt/hj5wfhHCW6pb26me6rdKShmsN
lOKfd9cvw+CVno+CwUl1AfqI4aYrqPdfIyXgFSPDDezJdkMqNpNINcYmNwe3PbZf
TGvfmbGso1sU50SL62YSTqvP2JHqsyDQY6fjjNDHQDeSYB/v9u6a3ADxJC3Juxk8
G4uq6pYRXngY5XQi7XZohA3q5edXQLT4A1Dg4BzhqZHTzGgqI2LqY78y/3TnAlsN
QgFU+KYuxgdipBpehn4K1nSQEqAzUglJ458MT8aSyxPVW2ylP3c8pwNZoc776C9o
VaOqoy16JzI4v9rnl5b8gXo7cpgXX6FhMdmulmxw0McFparsIoUYLPotIC71bdVm
wmhMCE9r11wfAMRQmKQiWzYqwvOAmPeTga0o6Q4qOpRuStNSWXW14dG2sXc50TlM
XkQWmD8P+Tl0DVKkiGuj9+dtr2DIFewbC//G3vM38Gu3SGvp54bLn/bX17S0PzzX
nbvg3AX3jXWERS051h3NghMjevwtLE3Inl2+Wc6kJlh3URYproBImfs7VwN8OQsw
tcFjvDzv6zSN3txWsyYiLKTwBh4QI1/honJ8FRwcQlfa9gPkuAOGoJ0ufR4iFR0d
yw188pjg5Fd5O5eZ/XVD/akGPBGGjY1hh1parSfFkiz8hJT6PbAZBChif4YGPXia
9Y0ARcCQPeXyDnIqYzXeVHUPfX5XSrim7jmKyPqYEI/x+HIkdI+zRqcFSXEuLW9H
JcOZuDO5tA/wct6K1vdoXCJLc1PgqA6C4EYqmrp2KYi2AfhEvscB471LywX1dfda
JV1h8BPfE2+PVyg51wmzg8ZuU3fo+zlZeUiLuxfGDe3PYahl74JMx8/Mroi+tjDj
iXTpkvaFgohCLb/hV/qPhv1ZZG0L6A5o4mpVgvgVIKv+4LPKPvgt4IEu7LJfBSZw
x9GtUFLxQm9zzYegQ+fGtMn90wefiF/fIxlQ5An/XQrkk5FebT+jNCp/dCChwLtr
ugtTMZk3gbkQE8WgZg+8K0aP7vkj+JKNqqJBZqjDSegHjsbr5cdMsz5IgVStAudF
uzuCQL7LpWNCTtHG+WyZTGvT/A6m2hzeHTzpDVTrAlmux05NiDBI9TwYGkDWOkJP
cR86DXCBnbb1cOojGdK+W6gl6uMme8ivDhhpygksUVfnqGLh70FvoluOCiSbOgET
FjyCqM0ZLspQcXzHMnnuAY4s4qRluXOVHjgOOUVs2lQXL6Mar2vBLTur2kxSnl8v
xaDhFI6DaK9Veo5XohZwoXu4v926Jdm10Zh8v8UibIKVthBFZcdgkaJrD/ub8EaH
ieP00VXHxcQcFaDjlRH2duejDkQtmxNqt2NdX89JfsERZ20u7VPOnaeL9gl1i93h
ekCi+CLrmqP5PS7FN/KbEhWscucRXnhSIRcUmy6JvOfGStNtgkva7DOwpJ0FRAnH
uMblIqmWm2biRRc2z8MlfJO2j0wJzVEolS24qs1thlrqdHHOXSZF0QShpD0l3Xx3
CvSZEkp0gH3xE5YxQfELlFngY7ZXxH22KpqDmO3CiLxR3UxbdMZiq6kEMt9qFtli
T+lY4ww9CxYUAcVcYSalqIVRcbAX9qEVKeJnMYRe1GpkfoSs0XuUnKTDVzBmNhYE
DdUHjRWhYN90z4wnUpL9NeSFLh/X2Kb8/pLBjaYzMKL0PX8NaW61jGNrjYWMd2tk
UyA07lc1h1zasyeoJ0fS+YpKWIMWr+T1MyYqB1xFhIE1a9SNV+iRYLABCfobC6Lk
i0y3d/GyYcJ8yKVB1rq+vlaowgrXa93MSi4po3IGqSXgLDxLJj/zKHlNGlmgpWun
fQGdGaLLN00Pic2DhhN6LUVgODhm9cCJrJ24OPu+BUn1sbHasP9Ct7+gYmD5EEsn
LfPICkGxjCtoF6AwWlCQdR04bxhgqYTMtP4Ief4qLj9hEVgnd7zWhxwO1pwNQdwB
Gl13BAb0n3ZDLiJvqtPnmkF8nMAvUwrfe+FYfHx6nE9C2h3AdiIyDbF4W9Gthfei
AOkrSPTzPMGyUF9ZLZsTPV0BC6a+OJJ6TISdbdx1T40HMTmYve7KyPYdfuzrZ0gn
+Vm1rw3Ft472w8eFwJUJXjrJX8Qeed7oyuBy73WsLz2UecFNOJPlhh9KMt1ZnQXr
fMIPMR9LptIfEylH7Fp3U1xWt1koKy5sJ8V31kZ03Lm69rN8ZfMLUAiLWdWJjIpU
FAMctPyLvjEXRNKttRSJjBrP2byWCSsPShpo2ozNejQkuRkFoOsaCD7XnlcRbheR
k2gR+5tCxbye45oF/osFfG6UVh97RKOw7ZjkiirAQOQ5YZd7EDXlbrFbfNTR7uJ1
EJYe789aF+cpStxiwBi/EkS6YE3hqibI5QsQfQT6iQQCLwSd87fN4F6g1ICkcyMY
WCMTmxSl9vPQp9Zj6lCBa4aDnIapOMshgrOmICVUe9ehtveEszX62s3hc23AYAZP
w4f4N5YV51ZzG1GpeOox3XA5VOf3qGT7unwgGSSB+wU+GgOI4DaBSqvNBJAGUYqM
3R+L/wlrq8X+Usj2Egl3Nj0WImT+me/dNCwNETvVis3ZAHXxHh42pEg1gxh9ecLT
r5YSNsoDMhz8aqzqqqdlqtk6OqCXYnow69XXS6O8Xopcxh6sXmgxeiraHvAKKPs/
2/gWOESVeqaDfHfBkprHo3fuN+ezUzmxBW8xxFK63RjjspCV8tsCvIH1hsh7FLWz
xzNg854m+nBDv1L9ERcQ5xhOD9JATD4zbOvRBWNI1+2VvHQ+YzG+9IHuSlXdd0oT
A4q80IuZIkzkKoiJQOF33MrWxdoRKJOIuUMf5oa+U8TzBFOyazM5chUpH/pHMZUW
H6N+aNmfpCUPCUFiQ7XZOnWBwGkrIVO2T/i+BcxD31FtPWHed2qzhBwSuwQGPn/0
qkWgLdc4eXhTE6mZIXZNLrmZ4uFkjbvoIDAuQnZHBrwfMl9MLct+cqHENRs3leEg
TuexfJ2MVnWyQmd5KAto0krfLMeTD1jXF5RaSoMPDtKpcX5bvtOenNZk8JZIz/pJ
0oLIotqm3LjKTz14UF9qoEEoLuH9hrttrSCiViPATGmvLf2XQ1PAGDCf6MNVDlQu
fIHzdFcY9AIJRxTv1pIlQb8gn/Q0Kqm/CZCXxejgIOQoYypsUt9xEf8ouv3V0Rb+
hpTnj3eNHHz3KIbmoY1xjz+tMCK3pBLUlMuxIN5F4ME8b4INfaLAAlmraroMjGoD
EUYqD/6j6Jpyc8aI4EQxCj36H1AdKaKw+q4WBySLLIqRVt9rRbggteFjvnnL71Xe
1l0bFmin5XbKxc1Tl41RVyTSttSpehdEmpQ+aAEixZewaF0wkqCfQQFOqtTF8xfC
Jbh8PFt7mv5assRLBO3XjDfxxjY8nYSVzKYc2s1wKwrulfyYUUi3PIoRKkF8+ImR
eWHi8DX0nzU3jciQPebDPJxnjqtmr6OEB9E7SWgHMOxpUTt1L2jTmhw0kp2qKlX5
DUj86ObCEtzmsxaShRMPQUciw571q8i3+MPQOxxSNUR52eJErI2nHUG2ahkulZHz
xH/F0nODq5o2TNnH2Qz1q5kHczGVRrSlDJpGOggQsB3U2hko7POZCKfVM2I8XjPq
q2Rt/tcxa6gy2oZFB5F5YcuU/mtMhB0palsCf+L1FmlR6Cz1B8hMmqAIoLgFOMui
bbASvIWyARMBz9nGJ/B1/ackmT+76RKcPCY7JtGjVkvbV7w1+HZLmLFxkUR10QiK
lXxs8aWn/TqKZvu+qJAB04ARL8ypJn/2yqt8qsAXiuhUxsnI9Mq+ExTZEb1QXt7C
tt1QUr2E/sRw4Mc4+mA/z0UcsgWiuXB1dydkUc0zLETsiO6jX+l0weCR1yud25Ef
lGuw8+qlH2u6Ws6Ylc/JKdAOiy7gc5rsZEyefhEmTTV068WJcadLYP376Kr17oSA
tdC6yGk0UK9ht2rZ4TY84NFVt6eg4qK/yLSQ5oxFvpf05pvTXdEx+XEsKjpRzuPU
QZN21jTmE5M7ybPH4AqBRvqSvVpWWj7FmwuLJFJoRsEFG2607OOW32/pMiJSe1Vw
/kk5kv67UQu5f5Y7zmvRMeXSKRvL7BUM4pc/dsAEEjT/lv47DKu5xaNm0zR7MVx1
TY3CIPneGEpnOfbmdmkddBkWClBjkIMsuzgtey0bofmvLpT/MjIpPvWxbFHymRzv
b22hTwYu3RxAQhK0ug0sj/tn7AOG87Xj7Oc6EJWPKlmO4nYPWWlGthjYQfqTtnpU
GvrtOb+LeaNiDAbnlW1M7HF6zeO62DPE1hK2S5cst5mLJOB1L5m0LmWnfbesuwyk
/uVHTyHlPYAHSSVy9vip3UtwTIINsmpIhnrVxi8wrVqAlcA45w0eKwHmIRx4bK/c
e0JZHNPh1KPZS2aX1B75ZEgH5/MXy+vpSd961PqCHKo9QAzfb/fFRQ2UWiPtTDT4
A/KE8D/2CIUJQSVrT2o4OgaPAQcom60MzEW0DeltVkSOMSqWkwvrOk/xdeDSZrtL
QL0gYpbfgRFD1eO9icG1VsjKGOrcxG2bIWIMnDr4sEcHS75PIYlPsPWATJXoX8hH
nxT3FGLE+jInQ7KPJJfUlhDxUCrHMN87/qNGzjYfnS5uQj/8NHC04Czi9/FoccB/
snnHaT4DKcJkBbO3p6vxrH7OK3nYcR0ekJTLJRgBEpvMI4hmcBMGgcwBCE2KGH66
K+CIzc+kWCASrJsU3V8YGQCG1dEyapwLruKlYEH/JBwLDQz5YIgKu3znkK9IUrIT
6eCPsl9S70FzcdOJhHEhjcp39UgeAzp8x7LMpeHHA+KHUas6iAgUi7sihlyjT7vM
SX1lhL7mI/KuNPchz84Ka+Yd86HzwdXHd1UaT4tBqR6cQcAb+4FlMkm4JeFc00iY
y9U4UjnK0YUBLMeuKObgL2/hqxbR1HWq+4ShqZLbIJJuvlG8FrL50GXgdyA/aM/H
WtbPYBTipn2LVwDF+1R+qg045erwWj7giTHHhtEZel3OihJhKB5nXT27sWc21yZp
vkfVu2ZvTNkxLaLgIwfWdq9kiiXC3CKT3yX4Ik0Xc/jmS0sf2rhQllGEysrS4T2n
Ih1p4mSO8Ck4uv4FvaKiY5cj/fHqIvBBCaW5J0+eWzj2pcg4xmrju+suwZaxhgAq
euuvUg6PREIj72USra4fbmDbhpnhjIKhSI4dVohDJ5T0MfhjocfETSrb+VJJQtmz
nlVtqva4Yp7zYGO4r9USnnV1BGAsP/wC5w35GmuKOTMMPZa71IxrGnW9nRFqxxFD
JMrjl+/MevlBPdjOPVBKxd//Th5DIjF3W13py36EmnPn+UKLDBdjcGUvunOB6pkt
RfhLmC5ORNM36ur1HR/iuS/DsvPhx7KheCGXrIZ8ic6Cb7uJzn7Dyw5ksGLiU3fN
zhSQJNn3r6D72Gg5Svm/sDGjfBh8LIfiEozT5VH20ezvR2sUosLtevwJc77xE2TD
1yF9Hk6XySOrH6L8dj5+WutQPS0AXnFu1FiBs7/3y/iZVJOsTTJlnxySc8gDmSt4
Zop34yB0EJlo8DxxLkop3c53JPNw5pEbTF1aFFFD/nLSlT6e/rMKrPkpcU0cIzFx
sarsUIByICf65u2v7mVlirDcGFLpbknKaAX66xyqz+5fkPz9FhIxrEd445xG9KfU
dAaBlRZ6sX1mWTzwVbtjlMH26nw12XjdH8adfqhoAGaS68oAO99SF01J42ZCOWGl
9vUCDjX4Vc63Q6r9nkcZm6U6A8gkWbFfgw7GKt2V58tMqMIrnKGP5QbB482chGB3
3J5THmyqdd43hbQNjfd4wBm99zsLhf3tuze5N6t/DCMqStL9/45vrysce6hLwnx8
pcsrQTxCnE4NxyKoCkFp4YmoX93XzVqQBg3ep1bR3k+BpUWIZAeSjrJH19WDLUj4
LrgMKdW4h3TbsauIeebkV/ovsqwjNzYt6nbomXhAeDB5GdVFrInWbA/dbkPKMjZh
jrZPazQYwirIMJVkuBFM5+N/rUm/bqJnACkY4meN0a0i5SNKE0Q2abgHq19Q6YB0
L/Iq+Ic5R76kOOEGZQ+YNcGI9kTW3Q10M59+j31hVo3i8slqERmTESbtBfBne8vJ
VAXk/u61lM7KWg1g9oI9UNrQlaeLqA10AKjLwjcEAkTruiHzC9W/vBxPLakkOUPZ
t/Ao64CMLwDsJZ9sJxanPkbhA4tIF1F2PzGoRn9goTKP4jxhafRbxbqJ7p5l9Z+A
5nHBa4vImdWo++Ypbmrm0yba4ZIdCMGzO/TYOm7RD0zn9UEr0tR8/mAkz1iL1HQJ
8p5gWQPjHpBAECh+8BQyQYqFxOQdqTYg6h4APK6pY3yN3bSrGZfCBOShhnhN2qqi
NDI/DCZikHyFoIrfm+I68BtPtXlbQquhSTQr4xfOsg++Mphke8X4mYag30PbUiZO
J5QUBwt3NNG9wihTHULrZjK2fuEV1q0uIvxVWW6Nmgoh1Ofuz5iaSKXocM0utzBo
NbG4p/Bea992BvogiBRynAzgnnk4KNUwOasmBnAsAJrzFOsj0OCNIp7yxRIIXX36
zOa9fgbT9SCA3xdvRRujV8X6cOb+wEigxyCLQiwohp/88k+97a8CC88E54DdurBP
h6yBqmQZkdBpGWHmkPjV+t0Uxz2zYa0/JOML4ZxB5DB3FKDg/4jgzZbgQpILy09i
eBG5vM8fnKVVdoc/tD/qSdXZjDeO3KeR67aZg1L3VzTKJmXK9ZHNlpI082lK1mcV
BLfe2IW/NcapSkw7aRP/mgjHzH5kiYgBnE0H563l3eYfaOOmOxH7bJxB2znCT4bt
EZ6A1saftMSImhCAyBUGdWq0lR5bjzi6KDmymcfXQronZvzaDmvmnp0o2Ltt9W/4
6w6P7yV6FCZbG0ggbwbq6/HksfyUE+QAluqjNl5I+bmevxNhVC7bhxvM7Bs8/Q8Q
e3Xd8KSDAShEcPoycEzUyt5Bb4u7QBDbj8AqOQQm1YMLHJIEIuWs5URZE2DS95XF
RVX3WCKVyK2cGjzi/xJxCOryJOS7T+oeiPZ1zpptuYeUxMRV7KZJF2ONDQDXcsyP
WojgmIlalksG7fgKIikmMQo8Ut/WcrNDz14mH4tNGqJ/UX6P/ZROJ7Lku1D788DU
rj4MC8+ZPu2KlSFdn9TZYPtmOwJxuoPni02OxayL463spv5IG/Mt2xRQwnKL03cY
Z3lDKmKnfOwx4SkEba7K57NzrY2gaqZjcSjb5KSoJ61mYocPqmHBt2tnA5X2IsN5
bXaf/GJZK1xHu2QUUnVicph5oagOxJk/M/88KdAOX9OhUrRuJVss6Md/0qh1HWZc
KjCCoBgoIzWo8vV8m2BeYznrYHpwAggbQI17X8qvYu9cRJh6DXRJkH1PoXS1ZkLD
0zrnlwn/NgrcOiv3yYHll7Wuef7mQrc1sUwevafyg9l+L+4hQ+xgMJcEXu0XfA1i
bYO+ll0VtRY7aD5cI2dR2zMr9aHfFESujAwYjdxQjsBnuA2UTEQDLbvEHx6QSoHF
GP34DU18IQJJZHGtOeKBylobRH7bLP0BCXBYMuu3b/DYYl+UZJ+NOSbVTUoA74Q+
pllGhmXfEFmo4Chtga1uE6IBpOUdLueFkEaNqU1QbcCaJzFPwQoqi37YODLGQELP
WQ5jOPpWg11P+/AEZ6n6spkdmQPXNRSepCUmzjsAmrOJgjb/zFJg/2OwD27kN9/B
cXYg10hAb3By2jqHOzbWa/xn+vtFsxEhPehWFs9PJ5lHfR59g4UqGrr7gMyGKZ5F
34TZPB9RgChVXcMYVQjugf3PK3wTZj9LhG9W6P06Fd0VT8qyEkQ+jMZ4iNA7n/IR
IermCPDAxGbp3k3TcFReQGduUPApp6hrh7Ltp3KQYVPOfnEUXQ+9mTVGjZGppdTN
wzN9ZGrHP1w/XMrNAcwTmRzP93NmZ7KCfM+SiNNyzblsJHE9KMfi8Qk6pBvGrkVu
JUsuHGqReVYJthiMWoGZw+PyqdvlhPHzFZdyOzcXsaN/mdqqilsbD1Vh+kSg0+Bc
om0NoS/C/qQlPJa1KtxZAQSFl+6bs4HH/vNIJsWQM9ugSo4Z87TyqrD/5cSKMLj0
A9JyA4tupdlKydSGvCpeU6BPhfOfecECVsZhN/dd6w6mlxndYonx4GiUI+z5hwfa
yg2S/pimHYG73pOd5S8VGGl6ZFwBi0zuq+iuAHBxbhRLKJSLVdr+wFXfxJTSOqZb
So8Fg7BF8zxsVfbUnav8u12aWVw9xdEPaOy4Yn+MPCS7KwKSpBKKasJIqU8TJ2ik
yR5JSvw0q8ymhT+WCQ4vncxhTHXn4TIcJ/iqsr2tiCVct0wIzQbsDia3OE4oHh+S
T3LVyzFifl5uEu3H6y3/Fn2IDGvukeA0Wpgkt/T8KmQ/QRlVSDCbyA0uIBQSe3Cc
R01izEeLEDzyTjmxiCosFpSRkaqkk2T3yaYVWvNXq9zx5wi25DDWilODbQhRZ3vo
O8ReGCWmABsPuz1RGnK/RVhClfNUre9Wammq5P8J8PgQPvqWGjnC5Sw5Qj10Y+Oa
L3K4vAj3YX9cDOyshqYzk2Jtf+2+nvdcd8j0d5O5rkWUZyGTLR2StlV1aKgQjBM3
oTDR1hZyYXlCafVxlYboUmxy98lnvK8CxKi40B2l8k/stKs1rNN5KvJyrE/jiyw3
+dejkPSOTQmBCFNK/mb7bspws/Vtg40sRxqpU8/qf2rTDR/cXzFLP6e3ZifLO+VM
gNdMJ8fkmIo8CJTwEsD+S2BkwqHnP2MXefZcyPA1ZQ+zYEFpZWK23tlZiTqHj9/D
mRhYGnglt7AOh4g4RQnbOs99wlKlwBlwqZSqhhSoHdn2hv//RvN1G7VQeaFMmB63
iS4tziqVgn4CNnD1KlOi4URnEb+pLlkpG2fU/BzgoVfMxiL8QsF8eJLjG9E1tPI/
l6llZTPQ1O9FNo8/QlbVHpMSHf4PT/3yN4HKtwzHhTp/JYeUHGRxtvskfgoYZjuk
tu0IkxUL3jXs0RKbaKLPSM526d6QP8cked0InM0vHX5QeHwJ9DEL70NBMz/aFqlC
GIkF5SUPkXsIpVOrOAz6sDXG8gL6KdrPH1VFYL4CWRjFRW6v/1KihQKGQPxdqA48
RgGA33mXClxp2vsan2jn5YJhL5dMB5FcrqIvZbdWrweBEAc32U9caU/hI1FXUThF
JCnvIDPLoTTmewrD634EKLGkHLBFBxlkWis+R5UaR/K8pz7DWXm64ApzrudKxRGj
CCS6iVTvqHkAwG7odn5ZbvYRJ4e6BDr4SihLpcl7sojSvAFjrghZnAFqbPtG4ipp
BDpO0pGmK/91XH5MxDa0MobQy6Jz9piAD7qnXC6KOEzl52F17LjHdtEfZFTlbsNy
GfYk8TslDMJ8dX7kEVfwuZ9XRG29gku3JVp8UHAIPjeGkWY45ew6KTwiFwSUXP4V
IuYK1Vegfk+NRsm1ySN0mdhEpdncUcPsqWPMs2hBqFH7SfjD8/zyIOyw5iEVWf0T
RdKA/emn6H0hfNOwvIwPxSnEulrzUeTzoG2vTMX13cAJflJYWOn3YBR8JSxukHbK
3uvgZz4b1cMs/uicaA93H7gXWvCfd3zGMQpvJOBskXtLrHXFJC7EO3X7a9PUa0gz
KhCAD8msiJ7dr7nz0orVHPVzZfZyh4LOevyavGZxWtxRNho4IMgt3/3h77TdSCEd
eT9cHlwkg7lA9+rMkSKcfoXeSBW432OF7mZTt8YAjSsExvc9Mjnp8hrjcRlxVW8o
mZ5G1O/3vPBmkWIdKTgNt7+jglEVFJewvfaZCqukGfRm0ND7O7gNnaFSa1DD2sTo
tBfhiXrNvCy5c+Dwp9SdfTNTUtSIgB+kXRWIvAZJ6laYHIjyqHJqdfhVZiGPJP+c
GpAFnOyISIkd9w9vyMSuwiSiVOA8GMllreTk8ygXQnsEr/uUqwzIyfiRwK0MJmLP
oCw3CA0iNSZ2E4CM8FHoFK0xhZgEMZkAsJi4fptlpYOHYVltYkYluCwsue3t7/tB
QNiSFkYP4Gcip5AzTvfJPp74zSFBjQiTYVG5vzVsmNw4jO8zrotjqlQhCV6nwKm2
Ip21LH9y27QRzffbkIqevFBAHFwn16Uv5mkg03j1KzwQ3rqm8vHCfXZPBBNTbboC
v6eSpuFJpczoz1VklSCUZiXy4X7yXp02T2aynYLJDUzS3cqt6goB6uTZ2tGYwS5M
zFwtDN3AQSluwvtZhvVyrOdiD9RXWsk2Dd5mWR5NmiMkqEFvEZUVaYasdxsxND32
50q+P2mDexCXq0iAp9Gn+JNfDW5OIhAR6rpfeXSKdPjKq70HI/GOU9eyZU9fzHgt
OFXL6NDAvWM5y9LqDyoMG5Be0/6hehNKtwzuNSxydDD1T/F0WO2zxXQu3yOGklvw
DJbym9wef067IYHnZSKDzZj6xBe7zNHIyv2eDHGRV9HP1w1bnI032dmmPuEc7dmD
BNg8othdKmr/4pBc0CivnS7fBMzCKt2yZwaKn8RhCoJfMFuTe+vCGzei4i6Xl+3l
rHH+e8nQazB0379moE0juX0AViIBS5WWszjoSmfwL2xqDeWYQ3Vn+fTG+kVMyl4q
LofgPjvp1oxkstsvd0g3WSa03ypWAyXHOShLkRTabW6QaAnmjpAx1KN1syrHpDLy
EcBfHMeD7FhhAzsp8IXEeFNJNWi3uYsVbG+xsbPGyPimb06NWltZpd0tIwGixwmP
yrSAtikEkf9VpbKNMqxvcx9pGBTx3MtLs6cmpxjckxiVfH5uh/wmHA0LHNbx0kch
CsTx1pPOiUc9e5Zn49QL59MoVAAdq9kknK4BXePUwtzwzt+lN1eC4iZDpnqt4HmI
+3zVxqBkIRJIZ42NGgknZX8VTK7GVDEmNnx9tVHbJHYFFRK0STPSFeGGk6uKvU/6
Fgf4ZObkHZJZyFszJbLv6SyRivyghNBPjhHmAFy2+DixzH0C4yBwbVJJUwK1nlFh
fDW0YzarvA4pzax8afDWyj6AKbCTvwk82okf1LD1+7PkggkXjeaaDGq/Rs0S/Xzg
PgAhW588sOhCRFHESoDM5CpN8Q7Bs0caFD05CFHinCTIk+jXA1PBYdCdh9/0ED9a
dXAxa+Z5YrtdtFiZbfuadqBUhkt6LVE/igLZUv5oQk9QXy3ScWv16YvW2Q+9MZB8
OLyTenwxITcJ7fpYLXInoZZ2NS7XXBeiAscywGgJh9pCHSjl1kzkUkl8kS6kkCLc
KQCwDkVSM2we5KS+CDbVRVDqpJEaAimLHuZJ/jyFOrDUWux6+CUIOxO+TUz0uPuK
nMMFARp+0wFBhz7831prdnlkJG2clW9xP7F5a++7lpVBCNlWBIyx37ds7y1a+9ka
usVSJ8uh91yKyyskKhYPKubItGTwMVDVnhCGwEAaNgFdDMvVEPpXX5m2Sw5PBIcW
vBCyM/2cUfGMBkjiw5j7Tn0dn1GPfP22DPKdoQzdkKrKLdYP/2yM1pRyGB12C5Nf
qYAOV9vOrd+lOHe3q+AfWWwfrjtmo3DemofJsVb2Na07ErBlPwPJcVNWZc2Z81Pf
Wf2IJIIKoCSXkhWd9JOaBiqHgJ1LBocuanrpActIx8aiGt+eHB/7vQfZU45smI5h
Zay1lnFFLOrEeJTh6TvIEu+Ag7VoALSa/vpuvXEVTuVQ3V77FIgVvN95lR1OxwIt
vWvurGiXq0Lcb7FAiFgixnc1kIeeUFOOyHTHB7QyxZy3eSkor9Ej34Rk3Z0dyy3b
yWnkyNq3Ci6U2tXj6lloNCIuREASXrwhnkYT3DAGFpzIKc//CFmbKmeSmfoAYkuV
hggWWXUJCiqWo8HIGE4i3gKdWqR/xMDMZ4D1GSLiVcx35tFNZNb/VnF/jXl7zpcB
byRzB3FZ6JdUk8Pe+6GvxN95QxJIlubNKKriBgzEPfsLphyqVg10xmSXexdrXoQl
Zod/i5dKLMfEcy2+mvh+VfjCTpcj9koB5H1kUzcPGljY7HuLArhFdycPEs9tB/Hu
SfY+78jIfiUobwNc9/VTJeI0KyV+aVt63enMiRHcRJZc/7O9Le0TKpqs958pmJY8
yVPYhkzVYpw1bOvqJWXhFgYemiFlQzms6sXhNVBAaUhKx72vPM8T+97CzW8uwG+F
pmdxVXS2HeTOCtpg+KMSueGz14F48Omjfnk1m5k00V4I0pLAYKLUK38KzH4m97bv
XGermVYMr3nKrSPzzZgJWjQxSB8J+8BM85KJAwWsaKTn80qJXmarfTJEmLg39XFI
SJVyk2UKyG8W0xTQaE8X3DkR9afUi3c3bL3Qwighh082nZc8VjLwbG0RutZlBy/b
M3iH2uAtaR9W9mtGSeVWkcjaA8Vw/yh2Ui1eXot7WPPdohUXXF8ts7tuMaHXVkVN
qV9m3kgTC+NxusI8cLFo3KzkcReDS2EAHbH0uR3cY4LetIo//hdk8NYxtHPh5rxi
dNcbSiML0gUAFETlOuQXrU+B6ShVSSyXyd2YfGqYVfvkYN11DGJXyrq3bhnZaQLf
zXYwn4fHLsDUtpIOu8NG0lIj5EnZdHe4QyVV1vU5hEGkTlJ0qjwvcAbKDj85+Pk4
z97oFjao3pKZDu9x8tEALtZnC7tsmAqQ01G/ZON1pW2ZCYz8Ptpjpj0050BhJ4Xm
FVVtvWCFLy09EbcZqHMNWC8j61V5fdsOoVZ21ia618NLhwpe6HDFYdQ/vJ0TZFhT
W/mZJYH1q6I/fORDjdQOcnFA6aLLcQ3qK4Cm7SQ20BzXv31Aro4P1s890qBrfuba
279GbLSmv91Z2WDTpEza3eRiBPkBD4qhCtG7KR1z8R91DaNpsGLt4pQktebH+02V
X9qNs2rDOOwQdJuAkPIdglbsAXl1PSayxYZX14F4cP4SmduIfQYQdnGjaAxtvstn
XqscdAvon2JVp+A7WmFpB/SBpwjiFnKV0XSaWKflDX3gb5LC/rQ5EaOGtCbKbYfv
JoJdNlQdDykGlptp86HP8ef3i9rui+4ve9zMsUgbOyKZtVGXSyDNmGcNHWKk314v
+VMROVuLnpnVK7jj0ezAHU7xRNaUfPDSc6xJ8yKOfWq09mLHS/KZtrU8sMUD29nc
MAh2lVkItt2i7HeDRvLEvJmmGPJUNbLCFkwioQ4xUKUVl9fKTk9YDtoGOiu7nmNL
R1RphQ338Q5LVvBp/bUX2J6CZOGclMHnBm8eTVJi+cQPg15BgK875rhAIJ0y4hYa
MXQoIk353cTRbmSl595ssdI9UkL1yrtnVLhnuh774X1H7nftvarvPI3Mn7Njvvg/
9p0c5Yz1iVRvyUwzZGxvpQQyBYKfbYl8t9VfTdUDeb1mc/MC5RKBp4sweR0vZOgs
EgQ4i6c5XeC4RiFa5fry8VsIHkhhCSCy9vSYi/XCn98nEGl8rHgVsDqFnQ9hil6E
wY829oAEabBUSJZajwNBjWDWP+oI4i8Fh5mk1tuqzVP89iWnM77WV+GfXX6rzQ5j
hKYeApStC4L71ntuaatQhpVvs/bO0aycjdYQac+N3r2u+KGS+uo9/8tDo2jzG6gc
BZ6+MM13rJOvhUrZ5CWjsiHDTIrqbquGQvZTUMUEPdz7ldZsnx2fRwDTo3H6kOah
v+nUWMXk6QJB4Byp8RKwVwAs1i7IWocMunAnWSCmCcuEKDkEC8YvNjEojia9yeKa
1ZYZaw9nHGdKrqJSJIOCrYgW/m4bgPWeTr04gseRvRnYLXFNuXME4QbuUEXIzq3l
PYFPa3kK8m0eOSd4m/o6j7tOUL3qWHUvyA/ydJkDRyOW/7+QXDUJf1owZ/dy0Bz9
O72yXYqZf5yjV/NvF9AQTgcDF1fb0ykcwqEfDAOtB9KZ0wuY0XdGZ6qsNq0OBR9/
Hb1rn2KG6gxewTXDOfa9SrnC2dHlx8r9cr2fDxzBQHGs9cyv26Evjs+dwZirVwRM
HuQJIpVThRYNaeocpneFDcMYXk7+UNQ3/wzMc5zoJpoiT8+4CX2lO+TG5lDuZF3o
JwrDoLzKUhsZnltemS/al4hiJaltkWRT2EQCpJGRE+zt0jTsISUftg1n8DvZfwfa
NShBLmqpaLNwZuRW1BNBUpFElZygTYQVo0tF+1NhEevOChrlpqVx2p23hiKpAzMu
X1h/fsCXz0wNnJ7uqoLf3TIhPtxb7/BaE7Xx5sEGhNmlYtFcEog51AI+BlqcfmiH
s+6UhTtEQTMv2W8fDnivRTTj8caoz6oPrkUw+0vVYlqNsIhkM+Yg8pK9Ly7nAChz
hLqYw95ZKENVhZ6NLVL6GHMLdEZFM9qdsVRZVVXLIVgkMvUzQtAZ8dHykILXG3Hg
1HXqI435IPjsJHHPdpYQpTNS1HGMGSwG8d8InX1WwcBerkkcpzPPFrEtXv4qGhoY
tHfoRM4vHqz2U9CLRLLnigBAp7C4B9qtyN/4vZZqdHlezkg4ij4gcFrwha4zXIuN
FYQ560rOZPO4t8/BvjGYpknt7+Zb2I7zEp4abZiU1gloAtvrKT4hYxTtpB4Spwia
g/qDScr6+OeuYpxNR6dXm9m+dr3gFccPsIEVaKsY++e2Aop3Zm1uPSFvT0/9QZQz
wd9bU2SNGEGrTCvZ2P7c6EB49lUXOo+N+02AOsyTws3qmr13sX/HL4aMLK//EKz0
hFgM8NQSXODFVIQRxbCR6MTl9d1ES5Lfj7tbuKhXoitzV27SURd09JIQqSLI2Gao
U/O0BZE/YaHnOwGIxbBd4UOzA1nR/08XtRJ0lttr7diOxRBpVrz/k7gL0CY8lgCD
hiSwuRObcQYgpC+k5xhV3n+a08tIgLYsnLIOg3/hUCbRgKviC1sQcX61FKoxrtYe
hjTGej0U2SN+bYcQ0LG+LHrrzEHv9G8QDD6BuFL8rAD/MahJIlnvcDlC1YqMdWRx
Iu5BlqcUoFDT/X+tWzo6yIUNFVxt0B3q//UTZEoqn1bPBg5ORz/K4XJQqVKj70MR
HrSWXOccqHWsdhHUGeqjroE1goCi+ABMzApdqU87u04S5aGPaTPdUt51E5elQzfu
AhiQ4sXqhcJjsr5F8xELaqza3ze0X4AAcvAh6guU4msL0HQtyOC5ZSQgYAyHGA7h
zOYkcUe0Pmb7cxwLNUcTMgTf3Q5ZGWb85deVQNDUTgevOe4wU0R/rf9t1EmiDJCP
9gB4VXAGwAoSKjrmATe+mYmAG1gkcjBju5V0HRLg3OEBMu66iy6zFB1Wx2vqXaFa
BMXdTcdq512oGvFx1b+Qikqry7A+MxZZwj1lRSNpBeL28DGcaWOvHhaRW0HcWchQ
8Z7V//mfxav+IpSUw3WtAQ4rKFYWqHyBiJ7hYIbxUUZ4IJAoWeaq+BfN6cgb+XMz
ll6qAbVipQgdbMYPtLs2lanlErLTQyoYCXKOh52Nsk+vMYPV0Tjdo4ZoOzaDedKu
P7pjwg8n/JqyxecoRUTTTV/Aa6nzSKj+QXrQnYgiZx2Xi24dWZYNMzssTPpHbT8F
dRXibm71dGxRRHa1gcb0BMugPe07mN3aZMHHwp1gn6krM2/c45LUevGu9GLgr25A
4Ch0pzzo/Fkm4LGFKCCFM9Y3aob78tmtkB094tKzH4rw5pA2G9JkMlsTg5GsCli+
2QGGLfZTWuXPj+mz7ngMaa/JeyAjsGRuoYnjNSk0AEwKoOuSO53cBDU7jmqQhlUi
V8UmWU8gU7NHFUMZgeAaLL7ULk+2nAnpibgxvaMgoHOm2s3WJBu+2u/medX/E+I4
HQ/Lfn3gblf4zmCwzlDlVZ4ELi7ue1hxRqaQQiwlQYCXBxTujxBCa7HRcCe2sPS/
Rz6jcMPPr1cOzJk2yIa8cHu1Q+qj122UWUdbnzwwd0WFK8rFBBjp/4IBPAN/Kurt
/XYf/xnNOXGgEahZNaw9i7+Rl0YfRjWreY+f2JS4s7GQDboSHkbG373Ipv5W3Kwg
tnRc5z+MlqChYjLT7xYvPCOCpSB5QqRJoUlseyEYdLwt6mY89yc7NjHS4oWNtxEG
BnJY9zoBXT4EnMuugpB3yT2PLGKMVdh9PlELXdR5Rb/sG0ttyl7AfmJK7Plo98x8
ly4yOueo8TuNLvz/qsC4zTsWaI//FADiNxW4sm8XzkyNN4OSNXEKubI908Y7U7V8
pbzRJzt7Y0zenqWUS9MbX3gunJO+FSWtBEKJqTCAt6ACFtwF7xHLegVKN1Ncz8T0
PC0Qs2CmCvuwaAs8jEt8KDqsqTLQG5mYO+IQCGqwtYWlpq/MJJPFVBkFmQOmNRX/
64CfrrDciuQghsNxKNnzjzoulXIskCuwhMOZ9Eh2sBYSsV9vk769eRrYoJUlD3Cj
IrLRn4Xx3CHcZSXTNSzVrw==
`pragma protect end_protected
