// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:26 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WGiai2DYK01aTVoqH3fI/t633x45tKSy9Pdy4RzlY5minzZfHyRfCcjaU56j+OXA
vYNeAUGen2fOHukPm0ylhe/2sA4SZge9s34mpELhJLRLzkshNQacCg74hbR+OjHs
3KXab3+owiMQTKLatzXK8SbHqBsMFRREY0agAyDPYX0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
4DDP884KACCRg1ziXjnEfpTjU7Zb3vjoIMzFhDhfFNNQuIXQ+onnI8MatapWGEx3
qYEsIkWHPBPyMw/P1Vf60Dph1MDCPwY6sZ9YavNe7BYVCxKpwY/hrkAk975Ywqjc
d+WPARHkcknByI/fsVvvVBfVV808n0fzJi3TIgmSJfI868zkCL9blFaM9jUi7+s+
OCFi099XUL9fGKrRYzgeEKnKpayIl8CUUAleU2cyVF8edxOM3WnQsAwgm1XDd0bV
22IsXOoyu1855Fl+jezL5hAx0xXMPyfMVH7iEWjuJMXLqLVHRy7Tsn32cJ5NaWDE
Md7hC9gYsyaUGzxuPKo5ITJeFO8Pl9Qvndt7qjvBWGmqszoOz+Vtb6hEMPH6CAxh
b/9duMkHsjEHsS0EU4a0laAcXi1Cbgp5zDKEbodlUqr2YXNxjWs0o8VCJK8sGH2B
MtFxsyvZboYW2DBveeSDuGZVXYSM3FUO8Xq2mgS3UqFvohvAUSP011U8S29wuJvK
UHgCmXhXS8CbuGQ2NM+yWWwFBqrjy8Wuv0g/s14c6VkBm6GltqSZzXbDlP+B2dni
JjdZlxjhUkfy4ms7TgT2bJtpPamcAmdgqckpYxgt3kxnuaVO5Lz7rxpQ1z4Okawm
3G+Z6Wywf9ITK3dip4HY1iLuhTJ+nNIku5jSNRkeQEGr2BXh5uR+e7Px9ftMnnvR
S7qK8h3ui5bAh88c0N7jEK6J7w1DTfSkY+gLsKL7Em6riF/q4HQgC1XVQdbj3CQ5
Q5Jq+gMcepwPdMgSaetxz255oUYtCfGF/TsV72f2WOnkA/5Ji2ujVU2LP1/VUil4
CNWZ5hwvHproF8DwMSiMkCR5rhfMd7QvgKXmvBsNccmVLgfw5ISCIdzeB7doBtnX
xr6hr4E9NVVUIwPXPvEWNZZjmC0BfIxDbqgql6Mst6c4dfold4HFYL+asExhfomd
mJT5P4F/4axyLLRKPA2GO/8JWdGcF+jj1wBDJa672SYlHVYwL71NidqfaIPMq6Ch
0tCxK85Mk19DcUTgrrvGfwV0NjBn0a8NUHyFLYvG4LZgN6N/ax1C+ZVlEvmdzMk/
zhx/TrFkvKuyYC6n+x5QM/4z+dZUFUHs6ghy0bQdFcMpmdqQf3c/M3bkEBowvIbZ
4NFzDObxs+0Rj5dfmJSV896kHSjQPI4SNRT4lHF5XMuXVkda0Ia+yP+KjJab5kwK
XtfPSl4Mv+epfKjzAHJEvmekNC9plENM+I+GXykBg1pJEzEz2o9uYSLj44zwTBmv
k8Cju08Izbq9g3dYfmbRcHRx+Qqin0O3evy9/sKZ+jtpNN1JbCJV79opTXy4FD4b
bwwEmYfs/e1UPnFzVt+ykEdUmepjmMjz9x/0X/HRjg+DB1nYvVk/2/87zAiLQ5tO
z8cQCkPpN/i+O5snGKM6zODVoPy12/YzjOnK2Mhp+lDiwrGS+vCEkb3SZ4hxB9T2
7NffYYJ3G/Maygs4I13iU4iiO8CjYi+dWe7h6xAZ3do5WJ3uFzQiRIMBpzjTZBns
2bdcSwHdDlYKR/zXZpZxwm34T6/ghpEXbtnAgH3VVf3e3TIuK3iDn7zf3jfeN/4q
BOS1jATZNBw0EUz+O4XomxKNfNgsIHRoMoCPTSByo1U6ED+ciEC9yHjvoNYGJ/SA
kZDShmxhVXtGnSpM36ZhFXvo/KpqG4s+xVKAtS/b32j1aJZILuEB4gHrxyzjeZrO
T9b56MmTEqFS3z590pyMCYW3coUu8NiG7NnWzNyQN7N2YMJ7p53cXMY2/86XjAQq
aX82HsQcnFgXxvbY0erDWQ7IHiMUOAcvhFr19FMjTydKKP/mZketdgvErmPmmIeF
lErJQRfNLJpmuAG1usGrpOj+clBDkgmk6UD5qUxoVj/5rSOQGIk9bNIM2g1Me8mu
57uS0rwVLKh+MSHeNEL1f0nVC+dDtPajHc0m6aXURpeAl0ZVpgL2ZtiTQmHe60Wx
25emyaxmGGPzayw/d7R31UbH4SejjhIPB/M/2GepKTsS9EWDIJ+EdtpLJcGNfC/U
chSSUKJ4rz2fh/rRmlvsUm/Nw33byUjQvOILErNa3xnESNxo1ejN8D0OrPLG63oS
NdnHiwB4FVYG2ZPhvbzWxHq74o/yKnzfCN7VDdEvvjsgkFU28Dyfw0rKcg/QPU1t
m8+dP83GQZdD2fRjQvLhdVMYrSJGeb3m2z1k3OzAWauCtXaT8LpbmF7lY1zClISu
XnQFhUk7Q3m7eDWb13mSZvMYyLzLhZeUDV+v9cBmJqUzhLhuP23cM0oo1W73m+Fs
wzfbAlxI5BcT7q7hnTqUH20DEwT6uWw4n5H2+4MHC+ERUhF7GO4XkNHwAygrit9I
C4JGR7GhLAuiMEMITewIKIyWjBSVfEzZjZYeNY+jxHLwqtUXTRP4vteNsN2J/Lh8
7sFAj1X/g5H9TO2hJxkZxopb3+chzVS2bMUYloSf/cLb3698Zi3dUI1xDT5dZ0c1
0o9gURGGkkmIxLM83mDXRycVAb9pp93yD+itLh53IqXv1MAer4RDIfOSLDBIvr4O
hQzd1hlvNbagUYAb1dQijW1lco/KVDFrfZcqvPcxaRLmSOszkkr/eY7kLnOCrtGt
fuFeUQG/lEkw3xzQbLULj3EaqFJounASmXaFGuaEMHXFMsTCeuTSq/GlETsjtbBM
Qw/rnp0gRJFOgyG5iGVW8mWMa4EI3feGjXa2PE1jbrb32oeIANIKnWYUIkUbIUbj
Trb36zU5zu0x958hml9LkIUHCiR9eqLIRhlXPzYIDb88S4v4a0/xnAsgIsfD66We
zn6+Mb1PL05SaAIYkLPIYy5zf7CKXGeWBsxWo30TvsDIa8OjxupDTVYJSLsZo+y3
k7eGQOQFb9BfzG0B/6Er6jboRzQ4ma+heqcTtBj48QQMeAJp6ib8CMit8LEr7r4s
b2/hULHFZN4QN5blxmv8LPCBn/EXI5acx8A1zQ2J9o471YdhQxL0JscyG3Mx1mSc
enxP0h9VJMs9NkhnTtqh6ZnUZiH79Z4O3AhFx5oLuNCoxVW8/TcDWpjo+dtOdNG4
RuaxRVOVaBFhHYtp4kzELdnBC84VDQA1P1ErzYOV69dZxfCiaFYXeJ7s/gtVpZYs
HZ0TZi+RDcqVarqhyp+CVEDG4Lbp1NH6mxklWO/fshkiCSkar3zoxJ5rxrs3Yrtz
99Lzr5/MtLl17fX3GivsPnPCoVqPZBjSH9gF1uMVupNReImR/9LxV+dZidgnKYAT
o1fnrUXOveBIODDKGv24/+sByUbKgL9YDR/QmonRrJvguDlfUmYU8TC9E5oM9N6Y
piE4UL2CAs9hdeLbBChjTHwBYxvRgJMO9m5rjxAaSR+rHaDpbzhm59hLyZdrnE+t
61DQ6GTS91yKoZnlSX6YLUzmvP2aLiARpvOqNByMZhA6qt4KooWW0HR0JDtimCb1
pLTfmCbyK9eWa7zsQXzeRVENPQBYOflpAlCkH+EuT7sY7qxpYff5ElXYyEtenoK+
jhtm+JhGTtG5Ik/mZzGqi2zyQwnOkL/pFbLi2L6U9Lt1ozIye2etgIxNKaKZmg4t
HviDOnEcB6R9X8TVtrB2H0b6uJiu9mhyCojz0d5Zy35FdOyi+UIbSMWj4Uawnmrw
DEhCcG690r9Vn4OWf5cfkItWK1aCiPCa2GFTwYTfLOSmv/rQOCewHqdV9Wmcr02n
DH6y2QQ+l5XlIG5d4H2pAiBPSgYvAoNuFNfAIgpayqyrAiHaRx1wE4sNeLpSxFfA
PI8HtAOu2IvZBiEYfwnrdSzUma2SkKHCzS9q0KfqEgbDng6gWmw4OOTU2RwSFw5M
luAIKEATDeNrVpcVPDYEV1JrFji/k+O5OuX7Q6uNpOetJ+nRjzjFCUf10EDSuZr8
XRGF9HJTXLPYaR2LcY7/1PVx3Uefi/uKnjpvS8wxp5M3XkZsLSgGE4WZq7lYJ2Tr
jo41EJN/yG+HQJT6CAtecLo1N2Jz4KmVXQNFf2kDyA8fF85HiyzSG2jLVLlLDOHh
aZY2qW8yGA72Ograt9wcN2lVCTXrKOqCWAIu2e4m/qg2bhmlJegKwo1eal+bC74/
xpmwOxNTloTssC7yYjzrkS8I+v3m7tmWuX0eoL+/ykv8lfcQwDHbot1FXXy0A+oy
EaTsEeXu4ZZoxMe9iL/kg3EEMAfvsX9YAbz05SPQVBTFzmsUGA7odPrT071+zy6G
lEXMRnVT7f65xr9A/pAe+vPOk812WYphfwbn7YVplhxdOjSGhbvh71ylxuuncQeR
Kxp2FFHiMQ4o1UOKo1buxMESafIMusgnMEZWlR7DZEb4S8DkB/jY+2wYhE1wC6XS
rmyUCYvM+52rH2ZWmmbsg6mSgvTINGr+oZQVFV/zLAcsvSHC3gtAjf57LLrwQu7C
kY8x/JBKHmoSj3mxj58yJv8YO7I4vNmG3hDbKXIdOBLEAwfqBcS2dG/wGkVgiCaG
CBorvOH3nWMITPOZegA8V/Rq+n5FF3LwhDISALfclGMbhWiPKby3x94OGLeeB2Zu
R5/zAGGcErCTLJsv8zbbmSif0ChCmMjI36K4J+rSgjQDaVyUjRHSpwDyo4K7bGed
7XBBvZKJjIZly+GLhEDZhp5sAHAsCn0YW4wRZ+T+PdCdVG68zt53NzROGacQeXLu
GPOB4fK4pyHfJkC1m6+zoGLv5ntsXzfO+NykrGueGNu/e75H7CCq3xH8WVNKNudO
eOpEGFEAAzxNpr+9HTnrUmOX0DB9voT6B/C1Hc5jKXIB5Gqi3FJAYy/deqLSguTJ
pFjvTQKuPfZ8/L0ydmxgT2Rv8gtshpYBzQG5y90Oe0qy48s/tmRSoowRcFZ/pnEC
jdt09mtQzSAfguRP89/4PQuU0/2iWPbQ76hh6LEbnhuUfJOysHUNMk/dOjszTaA5
Lkg+KN1aKQmlN7eTE7pgaejNnnW4Z5ikrnE56emp6HyLHiKZdLN+nqtzwvrxvnDO
31fs9ZMWnFfsIDEWx0P+9ClZVeYIQ0XpP1KAZ8XP3/xH4IPTKRVIZK1/ZxEUtvwt
RORJ+5aEyBjBHzHkM+luMUtgvBkl4wU6Dz/hmj+MGy4/Nai4YfOGoijuCRjKo4bd
p2rPSsVvqFa7W+DVqt0RIGdne5T8RTV/hS2le0pC8gEoOipWxN6J4YQg45EPToGm
/lDEBzOG6kWEvpDWdfCByVP8V4GC0GL8nU0YrAF10Iv3M59XiKf8S1T5KfSiY4Yn
AKwzU3Ntj/doHdQK1WIK7LGSCfWz0yqL1zEhKPer4aa0/bKACoRx6c0OkuiVZZYr
GFweV7enlOkgjanw7g5b+Q1DrykYQq7N/AiWeBJCpJvvgJ6lZtvvd37zRVKLetYa
h/g7ZfdZpiIRzxbtosSuu85gXgWNXch6aRMtxOKFfrQ3i8IIQI8K+FiYvZwGX4b9
9AKtwaaH9i6+UZXm1qCafMg4bwx5RF5a7CsMEJetd2X7Uo5gXO4FmkmPF7libGKM
c2HiWBvfZI145PnXRa33jtx35w6lyI3Rnc/GMoqeXeS7C5ahrxvV9XdS30dIVYva
XmBaGvp0z2GpA8yZnp3ygf+zINRMP5JH3w7YyWtazeapnj+DICVxcjYvoAbVJYs1
Fz/+8w8dMQ4xmF+HJHBVAvczqCUGpTujseGf+DtuKgAPosagQ7VVFHdX6m2tEqgW
sujP30KfLIf1sy5bf4y2kxY0VohbERki+DpWummsdwCsr4Ry0enHyp3MrbxZ4aJU
XNG+ePQSQoRs1H2nOhXRMjfc8t5G022m/RbH4+UfrbG1XPD7jLM7kpUW1PHdhYmW
psB72yxH7XQ04ZHdJiFMjieGvOunJ6Bruq/KJK4kxUpBKOPAKkxJmldGclDuANYw
AriOB5JzdGr+nTK5HqOLRFgDxwnInBcsU8fNmdz2SrweUwKWYbzQC4eTNZFA19fY
5Ar+a/wvQUdo6eY2gdM1xk0nBqKs2mILQRtzHX8rUhJCD3rUkYlo913NGI0AasE4
gf6Dv1JAyG3+QQmxvJVmvZiSU3sLKzhssjFMYLfNm8R+DdN2G2Y4bD4wy67jYbX9
/qoANoewsFuwcL4IYgod3+UufaiDo80EGuqnAA79wlkv/R3CUVUqw3vhcbVVl6jv
W34752CqogtVkMWe5Bk9krkeNZdQbd2TU74j48BqQeik8I2UL+ERWgW/dUWSSTYd
YUCJz0KYbyRpoImab7wVW02QloneFBiTicopBnY3SgclQfFmQvihoNI8u3Crpfhl
Hh9m1NaKPJp4flyNRnS2dYABK7dsXA5r6apK/h8RZgpxxNnD7yqEW/sWPPV44WdA
Ekhgtl6bquYTEomUMeHq8dj/VA345HAJMgryFjThrxtzQm80Rds9PvmWqKfeCSDx
HxcgbjY8okojpydIhb1RR4fuY5ljWa5/Out+8ByGP7ehD4oV75BYXUrP536SwekR
xEX1AvWOrfmXWzlEylBjZ0k900FM2SO7W0jAtxpZwSUACP6fcD/JHM1STsg7+oPu
dwzNqLZa/yRVw20139OOnB5UgqlvB7AOB+7AXABmL3PwLsirJwnJmhcazcNq3pqs
dayq77CS7Fo4nm0zs9wBSLIax9Py4oRMRynbKouRd/J1C/lLOQVXhFlye4NigMly
6QyMjGI5Q2CG69GcFy5uuj/R4r4zu0EdszhAAZUmWfxS5M4ejczFIQ7fo7/wGI9G
yXtVGg2HgvvQtrbul8ogS+aQjqm+D5V1GVwgV3V0PkmbfTUssuQAIVmlutQG5JeB
r6l8uldX8updoq9bOFrE0UnatZzHTDxP3IKzTKSLoqCoSNDn0tKTg3BSs9Baxz7S
9d5KYe8HOp7jvq9q6ztz8NDcxnAR+3KGmNL+m4V74RsWgcmx9/GqA+9v0DjAuKNk
N+FRtKoESDVNGV2g8FbR1LrEu29/GUNyU3zRUNkgcY8wDbG9K/ExWs8b4GoGQL/Y
qQAqTCgY7zFiEOzoV4tArhqd6cv1ReEkR/skll4ePYD85kmXBy+7LzQ7cOfddY/D
aFLIfSEBI9oiDTJ6IPOHwiTeMMv43noz9qsQR+CGUx1ZoK/dU7X9egBorkaglsUU
VKTXSXueOkmPX4DeUyQb6AXyutzUcVnE2hzditiBWHLyuGzsEehPzmKvMQpY7ksR
kY2rxeSHycg6uiX5mmuSSgE0rwU1VScfMbk64jhCEXQ/0MVAmz30tSzjoMcV3HgK
ouGRyOmdz3Sed+9nmvIbuC/WrGb65SjqI7FToUw3LOTKWO/cpqvcB36uBhkztvY7
OgF2E/zAjzwmG1pb/Z/VnzgUUaFGxwmWOOBbgtcq8liVMib4RmdWmG8oiSZOcq8E
GSdN7N1MmtkRCgOIAxPOsRl4ibaDKgEn5Zpv3sNXtw3Z6+X5rPDG6hHv1dH9zbu/
54HQqRCqTZC74CUI+Eoz4kG67r+hdB1jdH0fSFmWnECb/ll5P82a3eHnlB1Sdji5
hjIkUo6Fnw+RPRzl4Gf1gCQi8NZHtOCeDA5cZbnEuKX0mJvUtCwOtOwkrRHc2qrh
Nk049p2t1rYWWE/zhD2KxQhUd3duX1iOdBZjdaWt1YKKykOj2EU5d7tXDucpY5Qo
eX1dSqlTc7Qk5s0Qr0+b5RclbSoFWK1Xe8VB+FeIcOun+SR6pIc53FsQ4KpsXeaq
tX4isvHqPppm5ut3dMtFaJko302tkvy1AsTD/xkzTwUjQ596kS58Agyh/3H1ZwPO
xLuFvirj1qBk3lt8VIPhB3W17+hJx3MBaQv4pc8gi02t7LZNfzh+VypEUdHCKXgi
2euSt1zlPfAIiHBqbb1R/MLBNCSYymm0EcV3KDmDE0roohLJOsmkPKhIOgJCb/MU
eaa9qSkl/TH7JgqQEBjcmZavvtC+icxJdpYHJ/onXMhyHu4WNK13EN0IOG20nBV+
fLox4/leWyajRyK9NICa8HIeJSsyFv4Mx1Rx/a9/UgaO39CrDRxhRFmNiew4WkMW
Kpo2eRRfdcek3YnTcNcQfEGPPM2HQP0indtSapUXqNhd+lfF5WL3M6UsSRFbTjW9
cSRpO6PIZBtESxaGakZ/VCom/Exa/VnuH9ONWdqpW43ya4gl9Tm4cR7oOpx8gLEV
ZS8mmOveNKHma3l3hiDuHQnJ194VBwLMA8/dLLHTWN5HolnbclECIhH+RMvKCKIq
LoST71wMvYSxIdONzDGUta9s4Oktlc5dykLTztcIlDoEBDKVcDmbYAMMkaXBUg/W
y7ODGa+aRVnwVq4U1zjGdKBzQ4nSr1jixaIQxbR83TJSqL33VtU0rmrV98TBS+s3
G971P2wEou3NA12jYQcge8uretfVjRHSNYO39dbyk/V8APzPm0Z/sY7Fq95xrJDn
h3VuYgUVjImI9AYgfGCSEOFkuLaHxC7+O3ZLIgBS/UKikD8y+gkXVEpBOyzQ9d3w
5SIHNrfYay2xqsg+qrEYqrz9OCRdbSl/dfudIIRSMrb1OhbEBK4tI2nSG2xqdhuY
WqeZ2ZB8/ezkA3KcmJOK9tLrX7M1r/2LxnxoJdcRZWKy7E0STZSA/ALGNJ0niXA4
R0TmB2COXqYiVe6QzAuQ4du+2hP7B4/dFfWxD6yupFOU3TBgvZqdxZ9rQV9A2ndM
IYthjf2/G10lg5pv7usn4QR3bQTKC5rdZxm8TkQJ3isprM+j4ZWdaY39uyBzCjzY
hD9cwXwP4PQct3NmiqnVxb2gTMwscMkR6hXD02OMTh2APtwKOipTAHAows79cneO
RsXCX9pU1qzM0mEGmxdWrFMCuO4vkUoC7pi0JCwvsZEd20sss7oZjVZRGpDnz5M/
IEqjvAYdpbwg+4TiFUSQMCBAxvfPVPJRaD+AC7GOPEvUXYblmKetnctXfiU5uyTW
MJENDN+exiers8rP8sA4jEGMtdHtPjxQPklYcg7YvJmf/m96ZocP7fwVVY2yI08e
u2VoJxHL5niGDhWIdgAgPO0zVhyQN7PKJzTLAfKTmnA9ANChYAkCAX+sduAp9Qfu
PoyBE2dWz9N87v8asP702ZVtWQAa8g4IbNmyp387r2OqlZGp+mWBVaNSKgLBrxK6
dCsz59LkFwCC44IR3IIZQ7NMno8Z3FsbkUQxh2yT5Co9vU1yxzoyWK6Jd+QbluV6
wHXx/Loy6T5emN6I59qq0V2X2icDq91v52EOebJw8HXS8NmBkylW8ES5RhV2q0BD
FQoYPc+6XLBygkkI4lA3/TOa2YMUAAK27pVJgnBBF2ddsjZ7AhdUoQhuejkR3KW8
AzmxgbKpS0LV3QXqtlcqgNVrkEUrgJN//83oCjYICB3RgbXd6W5UKgWVTNi2oCXV
mRD5Du3UWerwrAn7aXThV+ka2x6+8aO6SrqvJMaY7TumGnO7oQmdsnq6VEkbvsYs
6+ybBdRA1hKrUbdNspbEJloyfZIgYpTur9bDA936TC1k25AQEd507YMfb0qdRhAg
2H5cfGSojlq9XYxUa2YguSuP9v8AuoCrlSOGOb4jPaRfTMQ2u/l23r/MsWayCTfY
fTCH66BEeuVFhoMDRxv2BtkazNJL76Xe2SfS5tnOm/JixCx4+DaOFtjYvglPYkny
N+IoPVX2ydoJXzXs2eFQnH8x9uYiZVAmL2d+bB4lpD0mkKYJelv6yP+tkGDW5FZ9
J3T01hW8exlg3en1Id+tpIV+sqItC9bSZp63eaaOuhO73RfEd6IWqr0VZvjb+byq
EESbmJ81ogjPtmDhYTMYB52KmZPlIEyd5jTYBmq0GAxAsoXbFQz8fEW5mUHbigtP
g/MxKgJBBZIROjlGxKa2fok63kA/5WTQoN1BaPn0ccEd84GVQkrQ9Y9AK+CbTFDd
0idraZt8rkf+S9KVY83qp9/Ro5RSsyzoOSaINBDJA1KaU5GAxPj5MqCucepR5dq2
IwXey9WJ4DmQXsfU15md7PGBMMwKKqt0MdVrExb7gijhZC8N8Wl0vOAhPVBvV1m7
UXODQ2GjHqSBdjLigaN+RagW+vpklplFpohoRtnq+KvwVUIo+Iuydn7GPPAou6VL
/IigBPnsv1iNJC3J4i71Rp1uzBCWYUsO7rLS0nphejY4IliPogXww1CaxUPLhPIs
jgReY1oIc6PUNxHniY069zggTJlNn9SwDH06JTbaRFVfsfEa3ljR+GeRtuoQGTkQ
8+wyyZLodPJ1acVTecsIrds61+vx0r8TuPfp8laoiXsqftqztqVHTxpxjtgQgycI
YN2dtQT99dW0wbw4mPXYAyxpfY7TKNqb5mbrwkAyLSD4zxRWtWbgoywXkpWe1y7v
MJJuDFU0XXMr1qPh2bGR5LeSrcS2VOKCBf0EpbxDqyF7s+r3MGAC0HzYBGmiYfUd
2qyHHnxD1+keK7DiGGKyZK2DcDEkMInw6hDhvgwedPCsXROGkB7XFkP6TUOPlRCk
0W2CW+MqHPCcPO0iY3kP3O8HccAOjqexaXZnO5L1ke0vB91sGWosinzrguG36MKs
ZKdbnvHckUibaI9L8/iwVTbMVmjjd2iRTXYMVuE9rAlcBBslkz2BPE3N8Hv2v9Du
rJeHB5QsbsxqiXQ4rKBoYjSFmfxhJZFKMZM2js/N2DQlvh0/dSeW4FzPn1RZnvXu
5nPuPVTWnNwW9s9See97noCwpGJZf5U9/7DuNUjKYleXWWahFZ9aWocvClgfvxKh
OaQKSzrBnJo6Wo/+tcfa/agOISbRsZ60ggwtNyAJebmgXeem5FYveJE4fFgFfXOs
b5TL+xoyPU7alIDxuuON9xj3IW7UYuM3u6DTJzu6wtUad1rEdmBY7IUIsZ//qd+6
u38/OHBj6VGUkiZNJdImf7u3WlBbGWHqBXGBojwgRLVcs9Kb+90oDoGp0/0Q6JhZ
13KwhkeRWm4k9dgHWO49yHxnNgvuvjGcMn551NE0CgVpuAWJNWaiyBzxBb1xVD0E
jC+MRse1egHB55+E4c7o4jbO0LJ8+HGt/V1crOfAQRihUpyJam3673ZhdOC+oclB
f+kvh5xh5KSO7OD8qMtVzQ==
`pragma protect end_protected
