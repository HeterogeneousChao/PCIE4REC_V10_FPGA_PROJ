// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:16 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nkA6qlbSFf/kG5LPz0McGNmGhmq8t65gqKlpkAwpJR1HEXSnl06HPl1rNY+3jLWg
53jxdC3vAtYm4A15rt42uckKA3E/GabONl+3a5VR4Xb6aty1WcGdnD0yF0W60JzA
BI0XjbLQzAWBPCTzxF1H1RI8J/0F4UuZ23sfC2BE2Jw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4416)
cxCiKh9A6VGAn/xF6mD8qxCSvbT4sOj5y1uCD92TeqUKeSpp1ziD/iqrP5OiNYdk
tSsDyAu2N4Efw2kEu8TKChh3eVs0WXKH2hHtmLiUOyh+/u/Tua4DEk2shWmDa1uO
BuFWkXp8tUzIqX4nnFb2Z7c59FtGTgRX2QPutmPAShU0Qi0E5MQq5mkF28uK1rWC
tXFEU6LYDd9zi3WovwHTL0xBdp3TfIFK9d7sB5jRp1Bn1cnxA0R7mkuK6KgcEvbg
H0Jv/ZUVSmcohS7Dgfw+H1Mwr8hHCBtYQRZEiiKTDUwC8TffYS7ePX0AOwMwAtnX
xVEURHZMxDS4+aRKt2I/czHk1r6X4TXH0b9XBCVP5MUQtXSWbscuH7J3mdKUVryA
DhUR/RPS/iKlyeFYBILTf2V0cbPlMfx1dqkrn4T942XUn96U6MuB2/mMi6thrPpE
IPBeTBiUJ/GpMbHOPDJdpDAjHCjP5ImLmXPSSN5U0hdtTC2VJn7VS8C5B31UfC1O
S5JxMxXir0goGrussw6fXDfPL03xKr2Hg8yKbJFuFmEv0wQHt+yhkeEh5WWuq4lm
wY77qGmJ1LT10qoEeJJiunlgBOpo6JZkm4c7r0nCEylChQQMf3KwmzXFoOnQPi32
/sQga+jQoiGyd4mCXRlIeft3GKl2b50Lt5U3y2W3ssclyW5zVqlBoenKVJQdNIRc
leFrB/CEG/gyukhW1yXzM5VIxUDB6Z6ifEcyD+1eFn5dcl4WL40YPhCoJBP6BJc0
a5XizTGk8LMkv1b6KbSJ+Oa5NvrUpgp7FxVgRTKgIvifrdJ+J/O7VC6TXbWqE8Ot
WUsukV826USzxOulpoTNaFmy5VJJpBCi9zauHBlhmsFYkV/sy73HONtPnoaMWRwp
zrL4ewMzlaUgzLzrBgAotmXQMiOrRlxjNN8flKipWqWTRVuNIoqnBW6EAoeCOhEg
pkz9o41G+byb1rW9i/iPWyZktkTbawgVAuntSQ0Hu2EFfZ+RWb4BCt2QdRHx4bUk
F91+PzUt5huRi8ble/PYolwptE2j3PLw/2kGdSNTCPtMFvYTHo0SWUHq4rkSaahp
Id559m9+Seefuz5nko+yqHYtsbSq8bmGsKzwF32BKlDRAMM3XWetn6/pFgVvs9Qj
zjZDyTs+MoIe2TKmE/6Cc9l0yxLkdIrEIkxBet5u3gKduw0NkCzYbILuS93LuhNL
Q3sLRL/M++Hs/iQ0O5SZERrvp7OHYcN4FwuZa9fg2UVriGB4ZHFo33ivM3LNrmdk
6R8xO4uUaliwobvrELhqcDQF4elD6IPqmTqc4JshyRjFJVbC2EduYnDSDreedl5H
nKcbZD9+8kcflNJFodZMd5PpYBC46dig45diWXPJIdezKECX0MzGd4XuWlweHozm
bOAxOnzFiOnm/RQ7ngIt7kZp4+Dwpv9o7i+XEpVkIGuVcg/cTT9bjySfySO6Hj1I
tjGsm8wp/kU26qtTh3BlMJ5DZY++NcW+egwacrAz8dVE/sDlWLPzoBTgF3P1aK1d
1legHLh0+Y8J2/Iid5FZFLQMwg/9kp555cOqjq9FbMm+1rTJG9BAb0Me2x/kYU9X
Wzf8omcSjabM3jAdKHItNwJ3M9hQmgya6quzuntTwhJROaFuhqXmF6kkyC+dkAaq
LjlRvK8f/DXGyWRlJOkdMJ1gbDSshRHIvMOEXoU+ywSdVq5lvIMlZuFc/QFuE97d
gw9HIIPr2PLaJZWDysHWFtLHATQEgcx2UOoQS2NK/wJZVQoMdiwSnCPOT/MYKWR/
5lVPnMmtivkolJz2UONIAPMWwB7/VJo8raqX+qxkL5iTp+sDswylEucebC2Hbrql
UlV2mFoehxDj3w0Z5+jdJMAk6oDbAnAcRajXJL6OKgSS6PYWrvpiewihicCr1kvl
RDOss7iHivLf5zXbjk6zrtrD235EOwptw/xtSBIh9duGeDwss03W/QX1Q3s67vpt
h8xWFusE8PECW6G0QyFGjvBUwEeHf+gZq6Cjf5Ox59LcQ5FEnHQ1lARPRaYXg9W2
fEaFD1pwkKOSvDxWw3LAg25BbjtMdiCsR9deA8j7uc/5mRLl3jJMutRE2ROmEOeN
JiK2/k+iXdnhK/zcWys1DWC6TGJnIhWZZKvKkGwahHa9b4agEe/QtXoFVEI+Is76
V+igkse3FkmFoPBJXJaMNcUQM4U5nsxhmn2YM/BVFQahaKmDv998sXLm9icl2XQk
2XvLbGNxE2gL36d6XsaWwYT3Seffh8s00T7Yl28Zw6WpOb6/JIGKC6UeNBSlWR2u
xbqO1LQqZzsI1sMBcwgtNtdfqD/ADnWmADj8BWMLUWEri9fR3bGJ8dA/Em5uh0ic
GKdlY5uxX0dvzwO4nM5XmM0MVn9zU/Fl8qHkuWV0PCB0s7kJk3tjw/8JxRVqD2wf
al/GZ4L3utnQbueRCulnzJiSU+96q1u5pre4xeAoLrE2IUw0T5acuN2TnEUXkICg
VdnvvTTqWJ8DTBolAFv1XS8Ox0RqaCLk+alHrVb+MsbuAhkw3xGj0Ecw+FtAqJ4B
R9Cf2NPk6g5B2AkDjBgo76D3gP2U7F3YnfgskwJYRVsBkP5+lbH/6okMTx1lK6OW
1PPF/thIQlvxpkDkCGjnMRwOWamilSq//eCxkgmlmyoj01+yy2Mu7oVMUMmgNwi1
lJyuSvJgcmuMjU5+wmLJ1aUvE4fmLaWkqOrf1+9GATAbm+lakAn91MRlNZpDOiAV
jblPWjnELDgDFaXJi5OC2KKuJ2i76OJ1gKoSTZscRpmRKoHCozeKyiRz3pe2Rcck
1vSPF3uz5uH1ba6Y2op+CYKguVSWNSzI6Nqn4s974E5uUmJHivBZHj4UT4WkcDxH
WbDAbihZq6L9JAfqvTPzNvFq59WASsLulyQVKE9NziRCDYApJ9BPy4YZUAEmGv4E
PeJTIYTXBxTe8fi07TR0hVLuTkQ0QeyyfaGXkTqYnY70cHBkCy6nDCODHpYJK1MI
WxONnEFL+5YoVdCO0Cofhj0uFFvztWIROjvbi9yclxpx7Q1KyMOKbANWb64j4RB4
M4eiTvjX+5F+WJA54KHHpLnjn1Ia2TaorVwbSVlXSbGW9wFpijJfNDXK7vgcgbqH
RHim7d7BpvOA04gJN4PtYdn+0hOq9XqlP7Ybdp9hI1DrWGzNb/Bz1XDmNHoMim/i
yEiBbUnDrsQn9kJh9xjLEQRl1V6AVtrk4PIyExyhC5EghurWiHf3BjhAwFEitZk1
WBVk8l54/STwhQeXAf37G5r3NmUL+lJIUlNpIn+/tbXN63EMlZUb7xgNL2iJsLtP
CaT4IfkxCqILPbh77cjMXAt4uL1INC0lVpta7iYE6TKWVZEj05sAZ68HCMcut+Qg
FYfNAqIABAphM/Qn4KqUmlQ5SZEcMPRi1xTwObAlhR7lolqMf5jG33bDgjFTIRaU
ZhavzQSVYV6M58cDzg93yBXrT7srJq2QNmhFT2nJ5LpHCgLzsm1rQ/wbfRpgewTM
G6Myz+SOihBWL+/tmhOhwlw0n4CUCzxPolfCbQhZlfUhTRDry6dk093QKm4x/fMg
AFp181jQ3KjYDEh2mdsLwg/MV+cQoD734HqyfU2zPAXVt2WInZP/ztehy949UK+P
VkZcELinHyzR6OpghjNR/lfoTXTU30IbLpPVnfegT5f8xfclmagEsAF7T6nEsUrY
PDaU23oo2pozUymqDw4+4fdFjF2isJlPsg+nw5GnKvibUON8XJRPCcrQuqB2uamh
f/qVYLyyWuYcXI1w7VE9hlmG7P93ZJYyD7W5C3oyKFGrmgS/QOgJngzR0NhzxHJf
xk0T/VXGcBmwH1cQRNchHkuZhEiTHJnZYfb5RKncqPEPpguiJ2ns84E+ZOelMFMo
ibENl5u8dL3Qahxwdt7DZb/uI5L2oLeqfdUBRTUMCeU9C4XRVUjh0+WfuNUc1ONx
vf2cXF7/gweX4n6WluHyk2K/oliv1LIVPMgnkAnxzyfPRZiLEkTEFzeEWHpaGZa9
MzhWgZzyxyzjoEbXLqJuaz14Gus75yDIdcYkch6ZGHrvdhP+ghqELe7iUKRHLRW4
JD03ZD3NrdJxWZy3xl2KiINIXjqNnL9UXJKMXe86l6UMixzWSnva1JQ6Da6VEXdB
TiWevJfGKkWsufji5kPipWaPY1JOJh8PRcgyYsvjXklHxdmN7UdJmvQEHVHBpkRn
ujkHE++STv4LoQiKnakTdTdR1arC39xUoiVjG0MNUXh4e/G09mQtMTECdB48rc5q
2CW/x2mLAES8bhv/KIz63GMo2js//5HdbesZ89gkacQPUt1MDRblLZwOzi7kqeqG
WUe7vCP/gxkLQd/27wfAw9SMT1QagK9HlvEEJ4b/jYtRDE+tRLvj8R4PdbNY1XFP
sqWd405ZOXGPRktPYTfaqLoJi+P0JaFGbzUKiRAckcNgiuxzw7joN3ihi2vi6YQC
ZevG1xppyVIcMMQ6EEhdrhPigXOT7Jl3KW7dGXYMDxB0WRtxK3K1642v9Z9vOACf
Niyz9bzpHU+bYc9TUqgUbik48NCYxtr2/TJ191+tLmW4ETbcre+g/F3Za7mqcaq3
gjnSRdTObmBtZvIJ9Gjjw4Qbv495z9FFKEnPScurnKmnC0mgqQucPgqNuiBBORhg
AJ60Us8tqsGKJW8LsrGKRnkACYznYkR3nEJhrd/YWug70ZDz3YPw+9N4Rtg5CZrz
v00L2sOfxEGwn1AfsyKDIYZ1NCaq/1vcd55WIqoRDEDTm0+1BNxeQMU3x7A6j6vp
LKBreMbeMbh58OHeV6J/tQfraAKwhhmeqQ9ysj1PIrKysIhR/n+/khiwGxon1gEi
b6HUobNzilNInzlh5f33IgkqBQ9/v1hQhMWfl/tqrX2K0unC6GFf9eij2I4NKRtP
F3nTGvnWLnLvheaVJppc/63HM4b071Tk7MPK1c9WkumEauQ+B/imTBzqgvW1bj5t
w3Uga+/jro1dj5+rggXc/iRKxtdl+g2nWIvizgfk4droOGDLmTtiEJEcBcuFAwD6
0bPMHVAeQ8w9gK4iazxGrgnuwGXv6MW43ABxhExsH4K5wdlgIYdQRKFRMEmhHeSx
L9DYnx9+c5Di8ZeO2e8W2+I2lBrDe2sD7/zylWngkeeGcom9wyMjwPLUkyGUCthC
Irs8wHSzjIpS6uVElFE9xPp6K3TcwEJNF+BSf+/EuNzaHIBNqY3QRKuQaQQl4bxG
TddTiTQ/0cBxnkygwVIaZEU8htiwuJbLkv90Z3xrg3lyz/dDWa2DpdSmbDbdfxks
HXC/k1ZSULrKmYlPe2pEGy1d00MbzlJgo0g5Pmei8DFv0aKPO4U/YGUyvwtAoXGS
eZBMK4PoLOyq57i+t5ECo4DoLYH70S5Z1ue7vac8du7Pgj/hn/c7rl10vgf8tQcf
qdNnSYSvMl08lZhE0ylAkz47f2UPlV1z0lKK7SbAvC1f+HTVktv7mJmjfrBm3yJj
2qTFHGRwCrNQyls96gVsix8zAljKHfFEORKsEGZMtm3zAI5jI0sfahiARe8t3X50
IDd5pD8CXs7EQHEmJxx0S2vvMTSiOgOxaSSfURA28UyDdg8INWoUiyYn53RyzHiQ
yQoJ3NErd5lPn1q3FJ1azYV7FuhWIG7SSaNBJNAml7jz997hWBlpoX2iAP6nQykL
HMcSm0l/VkXl0ow1wAPsSQM7CYDYP9lUvEqFeYh0hv0Wpj3uoIFB31y/d6AXgits
gFKoXfGAMTeFd78/bmDKenK9WXIx7D+VesfJw6Ku4gCwSx9bK9IIzwdd1SrGUnI7
u6iw7sv7R5lKlCz0HYY0D4pqaBnGD7gOfYdofRypC7AtvBlTlsQM2i+lXC9mKAHu
`pragma protect end_protected
