// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:19 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Lkwe8q7mlAtYdZ0xPX32L89YDakuSmpnfwlFjFBXPzaCZ2xQ7rVrGc7E5psf9c0W
Ke1KbqC6e+e/uy93JgUICClCjFZ4YFBVxQ9iztwxLDV4bBCFZyXMermt15RJ5lHk
g1kpeT0WfdPUd6OPYMPJ//u2HXD4jQBpZXVepL0hR7s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
O05WDvmyx88pJdqNlNTBYzsLTwad+DPg4q6tDsLeyea9eiDS7pRAwTF5U0sL6Xq4
75m3neZty5CozXRXaLaUXIzHE/M68+yNG5BwXHSzx7HAmwHFgS2fj1c7Fo9BWlm3
pZffwNq9Krvgb+jbYceRSvfaD9sRh9dUJAEG2OsWYQvKze1A1h89wKXOmPW5bl/k
fR2mwqlN/N5EtaFy8swzgflyyCYVLW8r9BTmTJnoKzXbJCKBkUBKStyTsd6MxoaU
XREbWe3jRexm2MQhmO7LZGdZRAZ4H5iCdPGOV6oBtRICoZ1mR9m7WRCVWkLh7VTc
YrEupRuGQoUzB6m6ZJ4v0gXZeW4i9Cd7J400f1/oexRNFk4PoQNckOdNipPNQC8i
hNP6zXtI3UBvORsVeeA8ZaQIAcCxQjxFsqmE9F4LOYBwgF/qHrjI6MOJH4dyPQt9
vRutvzdq5UODZF7a9te9KRPU8nec55R1y8Cdry8M9aGhyOR6fBpAeldFDXQ3J7fA
fDihAKlSWLHwbXwurLQYRiqF44Q3zMZxsFDrIsUIodHQ0rMfvI6ecJbbQEW4J6wd
dIBCbipCZB8g9xImC2QqsHho3iSVJWew5BQ/Mi5lhOjQ7PjCii8Sqg7d5VvMn5ko
hloD8PEZWAiogKq5DShC19UOvCGwnmCYrv0eqiUNW13S/Sg4Zdc1OLoTCB6j4meq
1ssiS/qoM9pOmIPCRlGsEvNUl0yo6lH4YuC/BJN0DF3DmsqbJnP0foMBWgw1bqWq
8o/i36+hdeIPfies/Agmu6eOaSetzN8DDH1jnLoVV3XvqmVlfOLms1jEdKyPxkbL
xaHH7vVMpAgNKVbMWAyPoMD8xtCHm6WUityG0S/AGVccKBGZndxpveW2IIDBlLD0
p3e84kPe7HuAsHg3tgPwHPTi0ve2z/ySpH0YioMDkwJ7AFtKxVkbwO/z2dF/UzW0
1k2EloVWvYr2nSGFD3gXgE7bWf893ga+KFYZ51ZdsTA5LxBMf6/HF5gOv8I+6Ye9
rl6B4VV3OBof3ZPsjdD3tkUybq0mlhk5uxbgUkT+Mc7ZFbLM3nWTpcaE8wkxgyFu
AyfYCCC3mHlocUYrM4nWqu32I96Y1k42jSx3BpPaJzE+HefrlNVN19w+fIKRb5K5
RkHRkIpRj2Qaj3zVUVbuLmUCTa5P4PoU5tYHT775Eas/Z326QvnuZhIBm7dHDXYU
uHEHQkbwyrdrBSIwbum3ntmN50CH1d6K7tYA1kWKZfn0R9sNF6LF2hpBG0CVcTo0
rQE4ZmnpjzfS+hmlI84QKSQvjDZgeniG5l1IXSdcSn4XvmFK0vqw8JgUuOBPPJK8
jVe6aCb3KLg/nYfchhgvWCiwATzWil4fOM4QdWc2Ie1SBb2sbaaGZJCCNl7mXimk
7KVj8/auTNuC42KX1JqRtpzQ/CyZoBE5uLSdLH/Mm9CpXaiGRXOVVXc61tCwp8bx
yYlFM558w1yWqX688uw9NhGfLsK7zvBjjTsFdyAl45Ye2KYlYp2xA555Zi41lryZ
yyu1EHVW629V30/8tFLfy6cyJmPTzjE546XAPnFGdEgIwifGQLdu9KoBdPtFAJs/
Tu0D+JOaUoPpxysZfoEqBSvWqC/Jn+/GwouspESVwUaYwaWxYSjD6qK2lvhVNs5h
E99s/xP4au5wFDexV0Qf3huLszvAp59AuDn3/za7fquZYSRZ3KIU4zp/x+yoseLp
CWsAiRdo90MkTReW943Bn864KuyjEkMYGxzFvbuInLxtTpK/Su8qdp4BnNhc0a+r
cgEbMBNpmE9goVqFOYgqg4YT9JI/a80gPA1MyVOtCE3PX2P+mmXvdczY66lbpfgF
X69jz0agzwqkg7tvZ6CNoObv24VDjI4zN7ZFtsh7KK7/+eIjP0HQjz8ibgiRX04C
vkKg36FBLhBLV9L6CVTj/OuEybzsgqsS/JGwVnqlpQMn2dPUG0yjvV2Zo2T4h2bs
jy1IzqRMtRLTL7426+jJzQa+YRlxjJCDH1UXh4y4VqbJsxMSUcnlhPtujZkMtINW
Xe2PEEEDl8Tj1sBa5KlqZU5ykanWqql0uba6p73A98sPdcBtp8d7vi6sZ6spZsyk
dFvD/MkLFqxsaw0d0qFHoN2u1JOmmDeZPtPFJIffs942ztLJhzkspEsnLTlUuyvg
4z/kAbMQBXDeLWR0QHpwE4Zew7I+w6NWXxB8vIvo8Vx0Wnje32HDTiueEvEEbsTQ
LpJJhYRAH/KmI9EQt/Pkpav4SvWVJLol3gpS1crmitl7dvZ1EaKUNfG/NxwgB+lv
f5n5cZqfBbh6beBYdon01sfUINfNji87vGsneG/AbRgh6cs4rSEjV+ODkK71WsyR
2it0ShhWtLYW/N3AOkwAThi3GVVRW7ZIxgx4dBB+BdHu2uEG8gz5BY6O9Mj3gih4
NA6ZH6iNrSUqfWlTJ9bv8QGNrOw4ZMaTjCAGCWpacpQLAYb79zIzwDnoMgKjEMev
YokLx3q5TIozY/CmF9XZ4e49WkDOvK9L6DjGBn1upcDLIONsdnsksqslNDaN3fql
r1r93jhLIe/7pw2ljmhOjECKlpKJqJuBKxLE0qJ580eVtxhfJ8xvYMGGn2e2LUWT
/Xnq/BmdPKvlMCbelZTdvLck6cyTN34SlRWOFBSWC1Z23X84G0kZ27+O9hyslRpc
pZL6oqqlXzofVrhEW2yL6SHBf/jlQbBkQGmo4WOGreMB3zLiNdRVEDjJ7X92kTZM
fqEvANZ5fe98Dzs9hCEy0GU4tWTluX9MiSF13yB7UqchURwFYsU2+h55cuTklYhJ
0ndq7DFzxFt83sIg2zHA0ZCB2f3M2GRM4HzTv6FsVAGXu+87ti8dJEFRhnEDd3Mc
ogkjiOBUtkstdPZ9FqJVWxAfOa9IKHfz2xryyqd3mvBSlnSLQzx8q8KsUjk4zfXP
y7996TglmlSP79/B/7/D/8htXWAohNn6l11IQPD7K5dcQmByJvfBm8qXgb+M8X1N
fjOTxtrZiKu+KkS6q1XmvalvrjlLqUs3yvg1bGWLrLOUox01r1PpHz98Al40c+bY
V6JG59whbE/tkXWq6kqUKFaKU0q6dxtztWfdDJkA9kZoGSGmv0y2k2o3t8S4Qwsi
ofIHMqkYjK7Q8FcGyrrolP3+j08jMJZ/mST5y3sqjSbGmh9FGWIWBVJ/MKT8VT8o
oQ1Tx35WJyyT1hNjggxJaePYE1QxdphqjnYN/l+ZWamAsITHSWK2h9AiZtJWf/Yx
B76YAlaiKIe0rwG45yS0ccuQg4ya1101QZrtn3ngNHiKrZV+aKdbqyLqydAR9Irh
6vBTcd+YIIuiQU1kqF6kQhmYsiCPDTWFHsWiV5NKW803+HNpswe9mkyrg+jp7LZV
eJy59NF61VDTscGYG6j0HPapRcjsw9lzF5DOQ/vr8ALEtDErXdvwqumAHwXOPeRL
7CL6d/d/sGwCOy+iRxghemAzw3coRgV/s2W/WTiRkjKdksOkbN/ITXjeDXFLG4EM
l/Tt4sMO8WkS4YjaT9jI/xkl/D0sXaS9iaJm80zOc4vnDzprETslY/0btJrr9ARu
FL871XlMCnv3mEdLsyNh/IpWnrHvCT/0vKiGTKzo3el6li6wMWefqTzNkfZ71ZLH
g7vPSGnEKBOqsElIM/nHTSLJgq4M0l+pFiMOE3HAdodqH3PewNTyTyHKMPujxSJd
yFuYDcEnEDBnu2k2pHU42y0SQfJQ9KWxYSwUx34Owo/TKgR5mUO03YuZ/8WyDHax
NvhnZXUBWJgh9N9BBlPKfqj7RK0uay5x0hAO+k2ODzX89M623m7BjsWaAgd7coOb
IEEXji+vUqkXVsugXjTS3q11DVauqgV6l6nnDSfTgQISf9YPlhXVLzYSftHjjHUk
ZEKHyKznaKpObWmbGzSWTVr0mDotjAcw1dWkGfVfBxVI7+s2rMSkr7Me+lXbvPDD
zYFn69nl6vFWXcOUKfqAvX04JiEoHGZlxQgV3mAiOBdRPZMGhy6XJyjjcwDEawbm
W9z3XQYeVW4RCADxIC1kM2vsIaBUc5ybxsgzitNHLnnp6kgrUACdzuhb/zuXKpdW
yHPRYS/j6XYaUF0rKGrlo8HyB2v90FGzkd7HQjVnNgdoCYeGarMfLH08J+P7hAsG
hOXUexKz4Bt9MVmmhOWCcTimdB1AjNLBMMkdqdKCHv9IY3UGDKULV1jGqfOHhkPq
pfaqL1aaBE60e8COSiAK/3Jrk04i7U73Chg2+YLQlMv9RxdmZLeTSwvEmhp88ohg
rkZSTxSjJEVpsumU52r/N7AxSyTH4pKX+r5//3rT631do7w1VHc3Qyw60mbnp/BM
5yms9f8oW7xnEC4P9GwOwb+VTpvjHZaSxH22A3N81U87cKkwlBqSyJ94iF8w01TR
bMm16AF7o9ztKSnPSGlUEC6+ZXQCg61S5lMPC96V16zpF8xEuN4aFCZf4WxQ/2Km
8stP4DT2L81/t/OHCPL100UvWGkEdfWY/muUROCeLEys4jQltErj8fFDze1GoCIp
Y//0jcxNvUGEhYN4nV6/Kvjx/NrLcDx/hL2xMuQkp8CJz0OIM9bBkBxio7mbbyNK
9sTWEfB7jQ4ETDGc+r7AxozytNT4P7GH+L0AvoGI/vMXDNEGYVJ+yg5cL6r3JxrS
xyY4ER+KpvdfYw5TIcZYqwZGpOAbJ30s9AWai/XJ3Nod8htvCFKD12+WBNsyIID8
XoCcGEcpMBjTrR4nAcwE8zC31rs6zjFGCmzC8wXPxd8nlfXG4eUhJ4ib12/M+pH5
pqB1ibhZrryt6edBCZ8VKmYloBb4yftOa9xOH6VOX1q3wgKrbfZTSZgoNPeMv+Bk
b1UytIxIgbbhEBZHsPQFfbx3DCSRDL2Km5UNzaFKveT7BtHANDltus3ZBlxfvcRs
n0SVspvY+Z2VgQTFTG4fbjg1fVy7maJqQqUvKj+otB+c3m0hhc+FO8KZwa5oo2Xm
FALMBBoDJBNHeQXlVhmpKDeYUsZClOSgwBFqtTNHGgOPWPAwKpl13gtfQpuPtxGt
6Id4AX3cl33L4r0Smj5HawHWpn4L6tvnJ0qqCqm4TmgRo+ouf95zyecVI1r/ChgJ
4AAOmhX6Ec7genCklhqLvdAFmiiZ6t0E8GDdTcyW3WzepCrUTzs1UgFU7DSV85LJ
20lke2V5qRDCUQKnXeS9I9dqvQ2rTYREo2Zhc9Nd15uPyl2H2cGgNuM8cnzBHvcu
6v29u7qO48sr02tEDnZKbl18e+sSKuInhqDfKNBrpRBPOQXlzUAAyqNJTBQMlM8X
eo5W1BNANTIEkSmumX2jnyUKmG44UlKfC2+4nru5LMd/aPyLUHntmryomwae0TWx
yPKkbzawOJNBuTmzQ7UUJO/DsiZHQyUm8bnfaR8TddDgkZ0CYZe5nWabV4uxXpR6
ZFTOFQuZeahhdl6XFelcx7pKtITYSBP+s0A8TVz5lFu0xrTfNU8LMqCXOC2Ydguq
ONWx8XRwsjk3njGSogpVI7lCt7FdnIJea2FYBwJXpN0a3KWCmHaxvOEq9J75Qrgj
T53Th83R1flnBUlf8+ppzNXQF4ciXPDhl3dkCSxFKUJpH2buNifMGaU5LuBmGi03
b7r4Mw1g381msu/wv8kKseVNyuMDsZO513rvZ9URMPxg/AUDSVetv5VV5kWfo11a
HeEnl9QCli5yWrYIlNMA/swIcNyDEGxewMMxNfT5P2oGr8PqzhU7H1LyYD8Ut/tu
whs8L1DS1c00DrJVu01vfZBqaf0nJL9HBG+pM3XhH24mPULUMuwc6OGzTKKuHZdS
xPUajyjyE2E5XsX0jNGhtOc4Wq7aJ+wuUXt+T63oJR59Ig9l4X7FR/fjZrF+yG11
+7V+ceIEulH8/uQB2ftlGMzQmiPp6UAr9Fo4lfXdqSBMgBjb1dJiASRpwJu6CsiW
6wRDijPQVHFmAXMa8ssYvez/Zg6Qfazeo+xbBku/I1oK1GWELaz7JOqPmTlzjDjr
+iU8vtbBIXdtOZVsUXXwBoRgzsbTyS44Mubo29CwGm5jHjEc9n8qPkD338HHVkUv
k6BH4INAQugm1WbcJHh1ytmdmbzQ5XBT9LFDMfEaqZ9HGlOVq6Alxaje6B/pAf4b
27Jho+1d/kLIpDMPgGyLD6uvc/KQ13UCnSD3hRHV53ZgQCbnrlsGYcSWD/GMEbGw
MOQN1U9wAYQ0fkKTaTYmWabo5iV4eSARft3rohTprRFOQL2X7WuIVDziVgDI55G/
tK1imT0dEVwMVIjgQ9xGXLP9UYz7W9wEsWQUgCKfTLsag5cTo72nTdossPdRq6pe
3rjoCPAGD7P4JM3Z445z80FMlALDw8i6/QRjTj6nuxBcSMXGTDDJtVwaXNpvNTmH
lou8r1gQAqeRJ54w91ZnI90JcAemREQtmMYqAAodLpnT/DoneN9LJsYLT75EdB1e
sCVQkyQnR7yO4bhM6QHAgegUkglPgM2NL2bVq1i49vO8DTKpfSt6TLZRdz6RMf7b
9eKztfdH2D/855cYij8JgunQFWHssi5Mf3TUUoBNTf+H1ck0oR14qUYXt00QP/AI
rqAuaMaSgB+cCzeCdOxW5wiafugZOFTJJIuhelsEKJ8SCRZhyI1b7O0L/5tNt62/
D7LNPcEmvr8PanlnKP6QAb/TG5YAuhbC1NgKJVfEW573NrBX/GYBG7Hd+IeetLsj
jOeB62SeZv4bzhMhodr0kW07x2ohkVeSvnQK7rVeHv5gUpYbuaWvjfI+FyxnYTN8
9wPOrcc+VmEC/cmVartdRPbrjMKLGkO96RC9ZWjk94kxCpziCpREHFEjJT4HNeMO
aRBfY43mmR5qvsWmAF6JtFo2BivObC+3llpF+zcJgtYL68Wmo+uAu8xLGghEDdvn
`pragma protect end_protected
