// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:26 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jKB2HVHW5iuN+IOE9YmC/zKOBW9GzKecwoRmh4wfFtpkoRiTJG3cqeVl9u+BSpD2
lxfXuutjMImaCAy/o3f7+1uT5APkDiDimocyJ2rfIgSUtgFTmiMwQTpRBRbBtYpi
zIKR6GHOSz7B5avCUFYveWeXegOk92CWj6N+MFt4z/Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16320)
wCSU4G9YUnu9u9lqy0lJp9bfrWlH5zaw++pIammtBdN/RKEMJtl66urHB/UMZcHA
DTxq3Mg+ws2ZDL0fU6t1A5BYwLy3lfhwa6jjsy+un7n/twrA0dA4RZsEpZDSJyBz
C2N3diC9pHeUdGIk5U3Ltf5JxAdHqdsg7+GzSDnSoRgNL5YUEHhe4gF0tbXOxYeC
0I14QhdKKZwyRHP2QWadBuCHF9e5n/kthTYKxBzXX9EeaKfefZlNekLwuw+E/G5l
K81lCFoGwRvxjTLfv0hURlHp6VKchSbNJ4TRKVnHgh1MUon/r7bCYv6tesubTYhg
cLtaBpvMu8hRv2siVgYaAHm8VAme8ekkQpPBlnxboVxivcEQEzGouGDeTCWMmE3t
xnL1lQ39AYGM29oM+u4UEjxx/nalZFA6+8CiWtsOVolGH/Umgp0ynQxqQ+I2QpIJ
kthyMVOQjghy9TsbITp8w/lR+bFHl3h8LRobhBE1m8qhEc5ozXHX75APZgRgZb72
hLJxglP2sQfrKxWdfqBY04g2YoDU20q2LEHsco/u6FFtalptLz63C/2BDuuwnj3g
F1+Tt+1gFLQ4RHORnxijYB+RuhihlLhT+7DPp3/cwYxrwbTcL+4PBZuAuI+TM00o
Q+DOsrYKWuTf3dOZz4bPZzUx2IlZ65qnRZ6XVrg4fIvXyyhGydIBpJLIz0duIsLy
21YO2kF/FeE+c6m7KVU3uwMPXMkJtl0Y8b2ncC2889i7klFEaHvmBm02oq0CwF2H
IuBLtcwyS9zT2nrk7GFTlIYaIu31znVMEzVcUwCIcqkIklhDpTd6unlQhHEl74sn
L2Effox+oS9GzVUfyT8kV941H/z78gdXWqUUSKrJik/KXQePhgAOdfSzvKt4YKRA
+OJudEHOD3b3Rvek8Dr2s3+9yRDc4FMKKeNKyaUGL76EVcvl+TsnKhOxXR+vivTO
x1awv5+D5hhO5kjrkysMiEnzin24ktOE7SvT513kQbKj02lcoRWNQ+7fM/oE+L8N
ybjfE6DU3qjT4gfouen8EAvThGBsJGK/1DnNRNFn4HhWtqU6cyJl7GPqSlyDdsdB
I+h78kUCqsEnOWoiB/2Yfus4ylaHPMRSn/LEzHqRa59Z3S26N7jp+4q3NQpiFsZd
WCUCD+yR+YOL1RNj3srkn5EFaWRzJK5RytKbrQ8WFd29Pprwj2nCiP/97fYa3F5b
+yEZesmmm1mUSWBP49rJ4/MHomPwjD2JilCcBdcXW6Ejgg7dhA1zvdBKJ3r6kcz3
9B0CpFvNPH5f9Sl+p+F4RW/sjtRmDKTs58YGpbWRBTP8Que32blkJ5K4+xgVY0gG
fZV0y94uDzBqM1dch3lWY/OkMu7o8aupLV8CTLxDaZ0qNHiz3EKRm/Ykl2d6vDX8
btbEDd0X08fpkPNseG5qpHy5zAkYBew1pUKrBhwBNtRU8rRTROsBGCvGpt2BjFpQ
xATps/NBcw2Q1Lxt6nxz4Jm8THPjGf/gDb+yV7PygOtpYR1n1rAUXfv6vGlM9lkb
KqPCBkvk/LFC1KsUNLnC3iVOPaczhknFKvJL0wCCCj+LU+hjbC3QFFsJq4T3fvm8
eeG5dTQV7laWr1lUbIQZAXE0N0TdYHHterHijDDIym5GVYX6Y3BLSepqqlm/pnS1
PL540ZyYPZ8uX566Al1NJsvgLF+Znhv7AlbjOSUEzBFtcFqQQLxRsMsKsfMZtGrW
bQ5j0jXswk2kaDy0CRvfIlvQAUAZ6QWzMn3htmi6rMGi89x7Lzi8Z/FCEG/aW2eZ
DUoDl3O3ue6SI3MoCWHeQCcQ+ia0VNKgvK89HqMeFIJ8hL+b6PTFGT6gsT6rTgd0
JsYhk5iLanVDuV42cYYXhJUdX9lU/t74ISR6c2s/NMrPvD3xK2sJGR83eqHqzRE/
p012XOMV4Sk5KfFwYp1HXYBpZR1ckeOKi5XysRlxGO76/tgezMe6qIcQZGQr/S78
+8vqfxF7VFntf1kbKuW/4JBv5uFntO5FTXs/16Tda3Xjf/hoJXa3CkwKXgfrZ9hU
VfcPWMZSG12SKBQc0kKw6T4+9cK6jQR7W/BcJvjCdaHxtXRguuLF7NVhIOtEY7oY
vH0Vhwe0n591ljhdBbVWBr6gTBou6+USCDACk1ATgXH1DVlEt4ZojCWsYBO0t44U
UuS/FEjYLs+1ClL1rInhiRJ4SkykpNtW39D4XW4uGkJan/d9A4mkcJCYDYGGLMGO
+vUmw2htsBfnTvrtGTGs4BhFCkx7uqO7itKp2ERjR90MqDx5nXisfvA8aMFDG+p1
Se27/+zIuJZd2i0LNhoent46psAyiyMgWq4pU03id68ml8Gt+jccLefYCFQHNgyF
e5HQWVufoaGifT3b0HOVtGAvc94veuGqoZ0In5hPUsSZMj1rt/gP4k6XlaqqHJkw
lUPlqVXVcb3bqYMhGjzHOMIpNUmLHaRHL+OkhB6ALP6ix7x3PrPh7z0MLYFEv4e3
tfvN7XzuzYls23SQFACN8+tKoGnXNrmzVvEcTrC9xpr52ZwP4H9j/elYSS0wfbhc
Z/y5Q6CMAD+wMkrhyLhm1KNEPovV7vBv+EUrI6xN8C77Jzfkw2tZlCTafjFSxIH7
rVc0Rf2cSgtAPQjzMpUICy8FiTEZD6hkqxKiBsBkWonrv2JtNRiiXSYl/ogzLSOt
RleX1OfBOhlnHjPqgGZwJzlMYAEGDzSiuJRMAMGFh0ISH+vLbv/0pCnh3MYfE5k0
iJdh283B3c9+OXeHmcYuVj4p5rSH4BF9UZRROTJ8SGsoyMipwTH/ONCYMCnONlVC
iK8Rf6/mzmEw55p8kF11vMazwnX7WzU/9I+4giB1NGEQVW0XLcc0mPhqiwOHIM3y
5LEZnsyhxlKR9ai7btoYD72up1eigwxqD489ywj44qgZ89F+6Ebg3BCdtrdsSMRy
BgolCQrT4fmoj9TU7B3qP56ArhwyrH5WlCBcrpDmca0plTIPf610Vwl40gRVxQiw
UGhH+dVdU2Nctv4jiVuTS8OC/xkdhugiEnj1Nt0vs+4uRzsygk57Cs7l4FcSOKrn
1Srrk2NDpOokCR4GT6pmJvQNXDlhMEq2QUFfRv2pt4bfX9MyF9x5Lq4oFu0GXB1L
AifOTkba5bDNJaTEOEYRYxR9Naa94g9zvW13SEGERQGwRTq3/mPMisUqrEc7eB/4
jMohaIIOwaAhvggVgLMoIfdlyp3PiS9RYod0sYi6BgpKgbLCuwphLs1PfT/Qz2lb
7rH/9Cn2zytj8riN1sM3fAdef6MuDkjt1tW5tsJcupDDUfmlW4J+ieWjv1JLXdMC
rF4UhGxbD8zY8Kr1YWcCUdgFJx9/1U2gxeba+QMjcIIanS5Glpz8pMwS8JixJThE
8h3bs62nKH8HxlvWipn38f8qAweMblnLTWaOgvZecajMDux5SXiUe2EfIvcrp0Ri
/zsfLdweqfIAGP1WO20wiWgsQV/G94ADf8WEDIp6KiJgs3vj3BGHeu62enrfIFCK
BKMhbJfZewHZu10TKNEg2jCJp4wya06kPnyfYNBJMUXZXe4qit+/kfvfaCitg4j+
RXOwtTZLvX0eg7SPUt7/8YgL+hUvHEXpNMFlk1Y2NKoPQYcrji00K+UzTP3G1AGe
kAtjCwd7xDCs7XI0TZj7/KY3tb2C0LUCy/Gdnns9q6Fr0Hs/RKeyBqqSsYBEpAG9
fDlxS0PxekZCLzZDL+8PujlvzLV3RWsst9XLDiJYwDovA/xh536oUHzk8HhE9Dt0
tU7WOZ+te6beaYinuKamL0wRHFsi+bgnaGqk4C4hqFPhMiWHD9u9dzPpDbur0gMH
akG3faQVjIrQB5Ht25B0ek0SFH6faCzWUi3dsvvwYy5CQ0UAUrCoO4tO2w3VY1eV
c4vfbwmMDC27+zhfoerbo/1OfU7VWkBiy3KBMiMEeD1SdImWpArmXpgMRHFCBjrg
4qYGx9Odfl0g37GSrcmLP+FD0QS6MbyZCqi6p6l1Amzrd2ktGtTDM2ZvhH3QOimM
I+wVKEM+8Nc0rtI0O1ooo/wy8HlF234OwJRHAuEzL7l4JjFBuAn00+YlSk8BHVRu
NOhe/dXjLyobKxxTPw2f0IO9578ivRwPGTxPx75G68c5rov3eSdMXzzH9VYT9EXb
u4+vP2K2EMhYgWpzhbF/ptrRCyxwcOO12AX2bs7tfnatygsd77VCijyqf0NrJgRp
RdUKoiaa7nPiFBgbkRUaDtkO9EwdyCyJuZWbRAtfRWw9yK967nzrVTGJRE2+OIQ1
iEAPZEJ6ldrsxp3yeLOKTvlRFg/kJsl74xFLosGr5pP/95l74pCSgxQ60jzAF/F1
FaqsMU5DcmG4K7ZJPzCKtwUGdLVsLkQf4tPKRVEtFqFKbzu16cYt/jJz9nAFGom5
cB0JZY4TDiZ/DrHxn0TMTuGRDPWx1Z40o3WbJbzCHj9DWtEFbBnEVNsPJrR0w2BI
QnT5Q9JQLTBy5x3t7+cSYfIGCsSO4ci6JokJI3BMvl+hSzXtFhO/s0/5DTgD8Eid
ZsWneS0Waeofct5MLlHnMEvX8hDsqAwjTnxGtXh+O8fi4Jn2GLJXNMD0fk84ysQG
LJNE12FcH7vhxM3TzcDxvYvDKeCvV11Sx/FPQrLG/3FwwL4+M8odoT4tOe4z9Saf
+10VwdJVNcrwtOAeIA7DbacjbtdcyYfJ/kLBmxyqxx6Oa2uU4/C8rQT7NTsYcLQQ
Qcwj6gEUTDZRlRO94znQPn8qqkrUPj1gHd2ffT5AF2MgrI8Gf3f1gdTZZkdcnHkY
77sRojhUTsEu4p1woKwSNSZDae/e3q/+33PPFpEwz6kxLe5gvRmgBLvx5mxGq/Fo
GEetlv/P0ycs+CjfjlMAhHtGF3hUt/N3MxTtD4oCRWbhu7aXJZN9Ajix3Z3i8jPw
uZP2DErLTybO2YQpshzYsZDjZLk6ZIo+HKDiNJa6LdhLSOOLCCMxdoimfBky+LH7
zeepps3bznRciBMvR5jRg/sR3gJ3XOlywUXmfMccll+GZGimS52H2XuVqJdGLAWQ
jOX4hLcrs9YUI2kEqWnrQmjNl4XK3GWCeZ0DqELCZNwFNO3unDkusHam4nVAZU2i
/wUwUYD33Afxpj0Tmo/zFGmFAIiIT1UNPvvsYnp5si6OeV/6y+Ao8et077KhOEZI
ccX4zR9rzkBIFHuKq8ohad/Shv6F7aH2F2TwEiJSpyZSNYLL1zZAJpck52CTC+kf
O92ufbeE9rsPUcSxM53/OEcJ95LRMl45iCkwaoRZ6slSb5gMbIsblMfKF0zIUygS
UWbE0C/8s84+Ww2TAJAWolaUUdNG2qho4j2lfhIecsuQpPjHlvqBWwhLZLtgv6j1
kH+mOHWIPbU2Lkoe1SfSuG3SzvpJb3jAw0nYKfD45GRW6dFr4B7bwCQDJr6E4IvD
ovs9GIQD3Ix7VLmmWJtWz3ytNPosOKNxSFiJhYxlcCNQzN4qNnPRG5GK6547TvtA
LKDNrBZknlM27cLHb2DUfKzIloZvzUzU7Hmt4SRRZZ/qCwK77dG6kQnySbgGLLee
OXcBYVqRo1t3QZ9qgLf87xpHBpOlmtt4xetzrYBgkUBvvskfRRtLWN1l9UyCNDxz
X2pJ731reQ8qDbM3oH2C/Np+XSTlUWY77XLXPrbxKmDAW6vRUhlcFIB2FOhczc1Z
Vr2KzLwCvGVS8MoAhAxJPN6ydJ+xQ1/A1Irrtewtw2ioJPxoYLarTiSIkb9jvZLW
7sC22Qhm5RfrrV2BhqmXzCCx1MAq6FnUuNAaCPhYTrqqAnNBva7thvzIj1MwKLcx
F2AXB1BuOVblaVqb1BMevEBzJ/JlojHYMzVJbL0hyoZfclWn5GvskgVSUGWRjZFz
Qftp2ARuQTPVDwWyteL9mp4qrw2omKD3bCOwF3mXzBn+e9XXmrh1AsrN5CqWanXv
OyBB7Mr0zIqAvdcPoQ4uAygv7qvsh23pfNLx42Q3pHxm0TrMEzEWjG/LR6ukewyN
lLZm9iAWy1esA03B6I+0oGDULed0mtY7zyEhWtYWDes8s/L8nyzcqxgcsVunn8jL
KXPqfaZAZbcTlVzUBDmQNy4Zuxb8WifoOGYKmNwsxD7ry9c+eIMdBqUSQwM8o9Nk
Re6aSlwQMA2A/Q2nEI2ZfKeYZwDHpIB+oqwqdl45WYhf3avkKHidV4jSgalF6cTA
Dx/rqw/92fzS8YJNpCo2jfjh1d40B92ize2jcqG2qJ9OVzaB88qtH2zFsAtq9ncQ
EFOL21+FH1kpnSIvuknmbaYkGOC/Rd39eBTyE0KMs/EH7xFpDeM/6lkXbtaZiR3f
iAdhHTdiylgtySke8OGPSmPHoQ/sqQHA8B25A3ZeGDA2fBxzVoQ62oOR9XpqtxOh
MzsgmWBTI9FKnPYYiYpLZ7HmD+4SBOT/ubTdYG5pygkmVZmdHWiwRT3UPYP+3B7z
qRLROcMl2BGqFdzubmdfNzSBqzSnCyBingdDKmOc5CH+WHLUMFTaXZ7ql3AtYaSi
FvfOEjvnOExxYwndhohVvUtrPR/ORM4IfKXcYEiQuTtf+A9ZKQYzd6Rb72bMQ4Lg
n+DyxF3MohdP5ojY5Y9o4y5r1rO6buK4fdeD0Nhj186OYA+zle9n9yVXs5O3p3Gc
QGrKLcyTtZnFO1vhKbKyIsxcCBjezqg7oYD5ss31dz/U8p8LoETnBkotgQEvGX4H
ucTNIInvOmBmDhX+n5wggKBcYoppKUuCLSUfUcN9D/LqhgqT541xWgdo/9OK3mFo
pRvnpkqORikeSufuGGvn10QddyM70llNqtfZNtXnIEaanGO6c9AT7Jc7MfUOLE9j
TzPlgO9/mVrX/lsGHbivfMELXWlv1mrxYdF4yI/CaBwKz/YpdhsrnICWgMtwuJal
2rLNDd3sSgL/ncc7GdGncTJkEMHAtkhp5qrtjkyswgawxFVHUkyv4Or2FztkZ+vH
lXDnTI3xsII19OUDRZZLS289D2i1p1kXCP74aLNpRFXIlFlbUZKaQ//aIVEouKPk
e17Woj1l6nU0z5D0RMt/xM6e0tON3nBL1TVcVZk0a8EF7UEK+JDaJesz+BUnbUql
o3cM3IHaT6WpyXqeViWiuhKkXYmqzlq3R4YWW6qrH2miEJYS0R1FOLnlls3cEXws
lSIV/CuQHwkE0bx8n6ZMlKEZC0s79+zYFO880IsUXYngNc3iBcW1SohgBvrHLIvn
d4QCBPs3pl6gRkwmU+X8X2AbgjcOmq+YQZ9lC1Vqlzn1PTYiH+OQrw+EPzFbhcyZ
h1UEafcWutyHVUuJlhanPm6qMpZ/Q2CU9l5a0ihwK1KdBP3LeHHR0qXRZtGtTiIz
X7rTq+9xhWu+Z8r/rZZVaWvpEu6LsNztKJUWOHBIJLlqwKwn68EK9mVY5Wk/4YSl
cQ7ogupvjKyhXbB5GtXt0tOOMs1kGR2Q70R2F1XbThq8uYddZL+UyjLG6oQ4KgCJ
AMALHvhazesmiNALSHtde817DEpT/fZFYL6xYYidosa7ZwJwlToKtpfybeTfVL8U
+pBgX1No1CPfRP2MVteUXLwx5sPHqtxWHdrRSi/IVAC/ajuP0JQIy++YnxcL6V1t
nHHDA1fHWFWQCi+R4LGEgrSrvUieCvO9H9CtMMfTBJr9qRDQWzv48T/GLPtuqNbI
M+d72lbaDGIQDphM+hyV3+hS7DWIFjAd4+qUEldIq40lhgHDzHnA8o2W5oCXsn1U
ZlSfYcDRKzJaxl03zuzLzsi+EyjZpVlbDdnsQHieNLCHk8TNMhNP5nnza/oDIV1b
WCzq6D3ulJ05kv4CCUbvvquVYLonHQeh35HhuPptLtTjo/6Og/AtXO1skqD6Qkcm
ng5m3gqeG+0SxD/VH+wOMxcE8pcyBQPD99ckIlma6rEj+y2a4BwX3TOvw6Ib34R3
nquL/Oph13wbzofl6CwQpNgVMwR1FjH+gune9KkFp30kSCIAxFFHZiUC1fII38X+
T6yWO4IlwWej+fWsvfgl515sgoNi4JaietFguYPe6S+lK/G4x69Rt0Cv9+9sDR0i
iBqxtz3sHyvQKfFVNo8T4v8okV88/I92nDouYR9f+xN3CPaUg0VBRd4FQZvfIosZ
KIx9ixc8SP8ZPIDJEoiUU3XdNUyAab5K6Af609TcOufXwZ/z57B0tQyQypqsCwm1
ENGmjppB57o42U5a7MfuN6MxbQq4N73YYtAvKeJX1i/vqLDdQcXaXee9uR/BgBHn
g44lBaJCUb86LXwgfpWRWeFTYhtDquYi+6QHNmUSZmErZvmN8Blzz6qhuHVqc0kj
XVhMGavsoj81l+mOKCUO6wsnDgCZHBMtRa1SuA65L4CH+LT2/20CWUfagYAqToXq
xIIIIaLnDRl3ah0JAugq28qU1FAsOXi9qot59ZGd6JNFSDLXM4Vj3XkjtMyNhD7U
7V+IvJT0R8ZOyzI7IU81efOuw/E4l0LxWy1y74tFlZo2mZkdoorfrsXAXat0RZI/
pvahDj1HZ5/OG5mLrYTX7PAslOwwTp8umTXpK/A8WXOqDN0V9k11PfzoNZiATtPF
aEiQcyPF0XGMztVAaqy0mvAy0YwlDEmZxZFnRsLi7uej2g68jUxlXuIXzZlArd7u
IkBmXTzKCXYpUMQ14D/FL1NGOMDLLqoyXXN128dnADkZPkNa8xuI1JDH/Ni6PL29
fAznZVDt8JiJmFITYUf46c8uXc6N6wu30Y36Y3gDAVLwqb2CfAbIK2yAMg85lHl6
B7D93zqGCM1EovLrJuhp1Nle/OWgIolwng44eiKdS3b0WFneSB3sDqquXvNVqs9g
eJLQKAnZnqW+NK2yfRphbc8mabP4J5MA7VIuBIaaGGmgoF6tf9MFDbGJ+sl8SkFH
4BWkFspW+e926SxEmcg2lLoc1mQ/CLINY0Je9wI1eVU7V99qL6XWdi16L34YxwCR
mg22uEt3TTZnSBRc9Zvu7UcOD2vWw1c4a4N5ENlZtSAX6JiB5/d/UpXmbFKVETzs
/cbZtW6MkF5lGTYbvhr58+GX7kzysUi/AYsdzr7+3Woz2hY/+VO1OILQIjJuUAT2
wERFYrQLJnaS7odzRRuHpI9j4RUJp8qGcDtsxzFrIzs75dS22TYBvrre8e5LRh3K
0YdufS1ZNCnCp8vb81XM6AqgfACzs1GCJ0lUos33gf4Qk0HvwHO7gytrCTQlvV1C
BxDWPzyc7l7VTO6RxwuOrhDoX4AQqaVofvPQLfKfrPc13Gz6AQzen9xYyP0+eb3e
APjjZpaHuuDzEe3gQWby+BTluXET9+SMVhqW+ePIv8h92/pNjSFynZ4NooSdbZY5
IN5o66YWnV2rCLZ6NV3CpXIh1iMJKA7NnOG6WgtOQcL5y/ZJbtB5m5RwPHrQx2k/
lqDk2Qj9O7Sir0m8p5t6NW2WHbKjzl06+0Pot/FJVY/Q66BNm65eALOdYJUK4pI7
qosztLW21dKSWZ+puzUjmmXGJ05BfZC3svkAs4B3GHSMXaJ+D30rBRY7sk3PCH0l
VI0BYS3nCK0aWSJt1W/y5YKqqD4oJOHgf4OVJhVXNzgvCkY5tjI+C6GzSaqkcw2e
jq5BECHVdWpHAjHTZX9Le+6ftx0t9BUYOnvewyAc1wvxSo1K8EYxTYhP8DV372TI
YYZIQSAPLGYWlUlCbvOp/+gpJQmZJ3F7InhJ8fB5FSn+R8LvFARdwAi7tk+NAzRR
fgDbqjnYsnHeyhVYLYx8E4NPZ2Iet84j/mvtNba53XQNdOtBxJwRm4Ez+MUJYd5i
HN7kaXAzbqV8uzRWOsVvQlWHV3o9GYlp/YFcU0kfSnWBABpJ21g19bwRF0rcANO5
Gb7AiPRgtNKcUXayZuVUpJq4VQzUgBIuy3dCd23X7mLeM3L1bTbtfYGk6Hl+CJOa
FteairdZnEBXF0eOH0avNKIUOvqORl+TFiWiyIj+Nie17gwF+SkDldLm/+SY7iz7
64znKymi/zyDwxUJRuzHe15DcIs2pvWhvoPtQukQBjqHzpvOIe+lv0l6x5r+kybh
AIuDNj5o/68fLvJ5gWGrCNlO+m8vtHfEnLutqkC8vAl7Qov4pUgQkFr1Y/v6+tGV
95AeLvKJpaHirG29FsQkr0oMW01r/9sQfnBeO8z4Jqdddn8g1hv0Y7irFFXv//pm
GCZ2qGr7ps5wpPIsLv35p7OP9iPijgBrhnIUf10x/iajJ5GKwYLkPiExyspIzDlq
P3lI3T/m9ZIMvp9PALyE142SrJopvMqk+DOmwy9QVDJS24++9VL2RGzSL9fFdHK2
9cMyxFgAIlL0KhcduDyb5zhhhjszbdgp5YItIlj+d/nv6HbbFL7hNK4uP+3k48gU
UNtuHpcWjS2/gSnl37JiZb0LL0UXWbQN3AVrjQItRUTasTcVGhGQJ6Ho+2greYKB
VdmZb3FtpvAvmE+u6rXmRQdxKI6Zthy6NxPBKxMtUVL5W1jmDkfWbuoQxaq46BzP
88qcDBlTB/QFO+NWKQb4OxvzPf2J1FI9lLhroFNTt0Mqaj95AgMMmIGcBuSyI0Vx
urGB3f3se6J+5U0TRn4wOl3Xrj20GJeiF7x3Wb7Ij32ygiENEL+w5s3CQW0GylDp
RJ5u09XYFekOA5JGsHLZjV+eSfDCt+lzOkR22qkQF0zb5qmFND7pzEWTY4bEviZ6
O2hkK2zmzgxFNuqBcY5qQ+M2NimEpBCxHMgmVxE12T4j/el1SC826nDK1VKXjKi8
8MgwcrYPG62Mp15fFT5te6MqJ6PWcmVn0rg4H+Lq4O53RYgAMHBycluFRufAyTZz
Zt1UuRWxMm0yldl5cWSscyUXzE7q4SuRUMELcr3IOZC1tzGal3Lkp3RlXO8+fQ9t
Tt7Cy3Kwx378G9uydHMaZe4uGlEiAIXko482EgWvTehQiEoUBCWOhBYgFjPAzVfP
AuKLOBauGXm7QUCbnfsnWy5jj79PUakzWE9ctiCFljZ9VmIMuPv03zJmMB29G8Vn
TK2LeiPqHDYUYXSJhVIwy/QmjuQ9t2YWh8sylwBxLSIy3GlySymudGUhA9qOLqcf
hPJ2Gj4YXMqAuZyUQ54WQ39TooDR5ny28ZHeB1eioxl1FWJYQoJLkQ8HsAGQ1nYc
BqGu4z7qxIW7WTFalXn2B4gZY+k8GTtRo89vPjBllMV2tcKCzGNiazc9eAU0CzYd
25PjH4LfwUhQtfL4vLOxdrZ/0q4x6CKzUR1Myd3GydnzU73HmxIILpHdcr7ko7LV
nesLDEYy7QjavoLqbPA+ds40lLISKiE4ptmKgHGkjklxXgPOdq4ZH6un6k591EJ1
qHOuiZpq+7sM2QkoOPvoIqknOfWXGN8QNhlwZM86UW8rkUxzeeM+1Yp6C1BcsdmT
tInvu1VumxCUfEbA8A9IQOXlOcRQRm/a0YKZ0tDM3r9q6gbqw2EqwezLsKio+2Cg
qixd5goi0RyD5WDYfrsoMkCe0WuU7C+r3RA6v8rNPQoQFbEL1lMu3nT2TLwjiJ8U
S95quhviJO+FLvxya/kZCYN8B4qNtqZlhRLzbbQsbtCxmBeRDxBOtEuYDcvKoyng
YrHllZtCPfNZs+eq0/6y5p1il3+Pap4s9S/8wDIwYRR/ULgDbvwywsroMcLikrdB
I5KD18t3GFVsI/RQtI1ITzYr5dQsELsaCe2Fx1Vl9zjwmbw07uVoqJZLE7gFmM+7
GuwZ82JJspv80Ze9gCyuzurhdWFSOMuIElHbpOI7mKD6pmfLQWCp9zDaThqlj3ZH
D6NWoKM0df0H1A0QHNcobn1e0eTVovgCOfRgnZ2M2zM32Kv28qllAUBEaI/TUR3l
yu66U2/wzDRRaij3euQKxRLFRC62cSxcScqtD9N06MZtiJZZ3N4pgso2dXJUermV
0upk6+KlYS7mAGXgUU+UNLjULq2MIDfpMVBKHTO0oMeVVTf9KztnX9FnEEAAkwOj
YJPnhmNVKFy3I5p7YxPy4EAAqHTK/RZ2UGQQrMkd4y1h0oUXTYvZwbjDr6W+Zwel
0fsPIr8p8UaZaROrAYJuT13QaCJaGWi5H+Ix1YUIJYvd+ZhGdvEOHlicEmPHS1JF
C12LOmqVZ5SEH1PJxgEV382LVuUJaDP0mde1nEGIkYdUN8fZ8OtG5HHFBuFKwg6/
kfaAhJ6tGOnsL9ai1dA9rf14mAXMgMhv/tUN8WYLF6RHVFLvEdcIHvfmgMYau8Mj
RPhRT26ISETz0Rg2JBHzdMZKHbt5f4OrA4mPDATcLbPacZRJiVrOT9TgtcqeoF2x
nFUJF8lzceOMtbCoJfCPz04z426iJO/tH6ENg/dK3rJjrLqdbFwrSMmk/32DtjgM
NA2u1cD1ukesK460PyUeKa1lwOiIicb1sraKeucg2dODxj4dPVE3E1Wc3206PEFv
SRVUigGBrijBGHhL92m6ipweTOh/tEBY+ycXzCmxsMKiHLnfyLGBneaWcT7r9pyq
ZI9QZG0CAa+7y6X227EAO1Lu22l2dZRxbE4UggSCZ4hYXD0sNVtLxWmgjwmbzEiB
iHvotJyve/gxNoybDdLZy/P/XAKNeaIUcUya1dbi5SO7R+3knhs+fsz9U9xVYGVi
p9q5XbFfmW9NCh1FGOneEnRk7ULqH5ApZXyPGwF085CnPbnFSlq8mX/BWkMAaZvn
k3JRCDxy9kciNlqNNSW5EE/bJU4h8I88TYwsQ6fJw+BpDV3YV1x61CHCbb+Ln3V7
A99oWldARuKcr7yYqeb7tHADq11WI4k+iBIYTpcztdvGczsy7nMKMKH8Z4gGOh4p
E8poDY0yJwxrvfyVpwVobsQp2Ggthvap2FiFsjrWqlHnmGI/Vmj5cFMj04vC5KKx
kEYD/QaYfjue7Uw7z1uQgM0J6ZhhrvyrBDL5grznOKJJTuefLxd3w1va8BXDrjwd
3q7NHAHH4BkLPjiijlr5U9QDyBOz+xAwJXtmzrD2LJ+2zgnNTdbMkUa0+bjdflar
NInAme8Aok9GFYBBtdlP4XEE4eNkz6ggk774vpDK4Z3e5095mnaci9x6U4nsxFvU
PKEeVPWF+2p0eT2A56QF9cwTS2PP+LUVJP8t3uxYh+7pLi1ZsKM2sXjuKwchTEYZ
a2X9A/C29J+xdCSNVaF+Kmgs1VnhDBbUQmOAIelVfOKoImglFX5FDSqLklpNtKMs
phpDyXJD9nAG1pYPlKy20luYiqLUczDg4TC//kmHBLrPuEHdlUbmDOqo4xqWbZKC
81ZbpFAWETFlHMHsPz4+m/T4BeEktlExxVfsugTmfNgQwM/zZKLzdiXSKDNrM91U
qxW0d1L5iEHxYgoWWVND3XrZQ5iuXVja2Ge2NKuAHSkcdwMy2FopyYXFWoqBWh3n
ivn5qfafYw0hV79p1XH9ucFBUFNCQtJj9U/ABXmv/tAnCba6wNtF8TIg0v3zXKYn
6ECOq8Lf9h27wMsvPYVDflr4E5bMAqZWOntBILHbJ5Z/eSZQ/ppfJFDB1r/F2GfD
Gin4LRHdk9zb05giw+jeO1d0aH1tzoCyh8s6lgtRLaR1u4e6WpakwgXrWzU/92rv
m1Z1zwjwJJI521JDhvpGmnAuTMVHl9lgMKAcRZO2kxnNprVNtsUjB8dpRKFb/LJP
Qm6lOumjzXtn66esnNAX1CEPEKq8+LuI0ZJqG6fIJ0lhTi8/uWbS/3PuKmEcAIXJ
YfXxMQ2RGVvwkkV0a+fB0k3WGLXz/5LntXy8FNHkQD1C2MOo1fHRZA2zc+MphGDo
L52C+Skv8hQfMze85mBqea+JKgXcnLlyY5EFPbuzqHDu2Y3iwmLw5f6TdIxsvoYF
g4g5FcoQn6VAZOdPL0Gd5tX4Q4AGbQl4Z4Pzcpcy6tIDPuTEFfm2egMtIJfEzDP6
AFdyJNqDjzKIpjMvEz9P5InvclcZ0EG4laZGEzAxWED5i81y1dXH/xM0R4SkQli9
K6ek9Pz5ecFPBJ+ZLHDjoLciwypSW4kRnUiBc1EDSyf8okTwPJYkfEVchdblXMUR
+UEAzU9X5jT9XdJ48JJRkM7FG/XPeZhw4tItz9AXdPWjcEUE+aDCQ1j6nwJzlJgL
YarNT0D3CVTXUP76aLQ3YNOsJZ9YXw2XDFcnU8L8CIs6QIpEPehgADVLDXidNKEC
Oa+r6rTqiD1MuNwFYFJ05qhhmjZ7Ppikg/EUuFFEWF9gmn+KGxyW6qVb092oYvKY
BDbsgQgmvRCeGio1MBxO5AX86WgIP+2NhqwUXXKp3sjFaMmtN7Geq4/L8Tj661+F
sD1YGPHc7+zmXYkblZmszQPJAPppEeXlaJFzXnYALJ9rXz5uf+WXUVeKIjFWtjaj
UGHGUSHmz+hRHTj7RQh9ivT/eVvt6ONpBnyBMLdTh3RyGvg1h0McnD5SxoDiZsBJ
V96HdU8bpiELfN3ywntwUbeIVTH+bH73CiuB5PbJIHLADAh51zG/VB1t2JmUSZ7q
nE3N8Ru47JELWSD4IXmbIHA3Z/xxOMFU4PylAXoarbvIQB5LbauR3C8ULdEaK5+N
V+ZSedAukZ9Dk4tqWWDm2ooevr5/SZyiufmLB345zGpOm+zOYvXgPptqlghoJwW+
as3hcZ+YE+5ejUkQCIbsWlCDhjKlQt2XNtLYa5PMdCM2ljMESUGl4BIQwED42WYU
ULtDM3WR5gBaV8VxGYiY8DQrYhq1qWZGFlXtB3S9VHXwdzXS2O34LdmbPQEyBzea
GzaG1QQ8SXWGJjQTR5InSEVQyxbMFK0GLz4692YmBophFNVAFP2mublY00OXVBmt
kZpG/K5Jfpb10BRgaJ6mXWcMaEuefJa6ZzRDx90q8HVW6dmuX5YkQhhwsBgKKRL2
ww9DMrEXp7T+ZLw8JytkbbrwChOeDNdNnXpDjn38r4C8wqmOfmSwoZLRJF+jbx9b
A9PFZAp8wLK9zdJtpGJrrP/vzn61gRXjB0nZUPZg3lPeSqZttB8vSw2PNBX6aul3
65NmiY0kr1GcR9kxV4u6XRNp/6lxounVnk5yt2J72VBdbMmk5gDKzzrYP+0ZANsr
+HgRga+p599sH7+SmjIk9zfpcVRnyuxs6v6k2P//eGnWO1Wem0CpEMYBL0PCqkE/
YXPWPNSin0TyNrrRcF0PROkj3YwdQCZKEKdgXVTUfK9O8YodyDr07gUAvDlj+UAp
xKIFD5ZInbvU8BFt3ITSmwp/GY8rvgfYwvZnguMugPwrIr/u2kt9lSvFn9fgWZO4
LONY/mgQG+gRcwwFgHh5Eddpo9GnJ22ze5slira2H5k/wEuu95hdJudhGzVjLldj
tf55PdsBSsmDlSYN6+3IRP+tXGcGect4e+cdN0pk1wzGK8cdjkg65KGRbrP4yASU
JhRM7EBbFzr94TA1MXMYPwrNkFniXIIznePy75SW/tlU7jyQ5HdlSExH86neEshc
TXqy8svJ43TZZvo7bfBYTTqAPvLBbcCNVq78p1wcZP0J8i5TQyTPrDB7CV6yLMmb
UgPa8dW9GfBoSMFj8cJDnRPIRsIc3C5teBFlvYcsLlbYj+eCgc/gqFZnBGEqCt04
+xMEy+5WjTeF8JUoHoJLy/csLTDvs+p/HWgqivMPx5PivPnPl+yJ4lo3QppNothf
FEdSpFudqGl96/Y+eMH3+SAryA/Wnt4l/Il6NQdV1tc70LO7jJKvtPY8NIqMqtQv
OGmyGSdJvRYE36+SPzLbeK9nRb20VHfJRNahzcD/LN6YZf9BZ2pcil9+r7gcfUw/
WXV7MHzJsVfCZkAGmGZbHJY6hVjJq0M0LtyvMiFLPp3SxJMs/RivM8uy61DU6Bx9
SZ4mNGuA38iuO1mkfi1WcxoN4YSedJ476L1FABnO0pydlBVVPwtZUMqIOS/gSEJH
5DW4Z0UFenWsi0BiK4ww6ZekOy/NqWTUJQPMCyjd5OLmRNS1H4A8fAsK+JI9oY6V
egx+3/Bg2ZvHjAczSH5Yc5qFxDeauVsS2pdavzhMyTnTfmc7IKPczmA9QcNtQ/w7
IfV5LSyVENkxWXi5bON9E/haFLxEYA24/ZBiqtBBtakYu9QuKRaTCcRuXMB7cVFH
tWug47fkGURwKfESI/jG4+jzZp+gswQP7OqDUvBwkMwDBFzYBaTbSx8oTfh/Qv/k
AZNN+t3BSsWLyEKvm4ccbtUyO6Y1v9qJu5JWoiExoEDtxU5JmS3WGPztLCHfgrql
KeRVwy7zsnk+Ek/rUpg/aRV8SVnQKhLB9Vl5zeMxOA1wkBBFe7W2b8YszNr6js9+
EruS5ZU/WQdEopwHp8a9UMFJ/dN/Zc0gCdfHWZ8qAbWS1+DtpxioA3HdHjlF9Lyw
1W2TVelh44ZPoyRPSL0mBjt78FGCJmD4xPAx1G45yIRcODNcBrLgiVQLSAj/2kBU
WZSRQyD2BcyjgpPla/TCbLYJYe/oA5lGvPBwNlZz9WjeU+eEJZT1AvVYu4JXoTgv
fkoRE6ZBEqc1D+M+NSMQ/p6kHVJsYbp3XGVXjjSwaxeSNh1panLHqv9dBmip9kCl
14lEtcolNTsev/bXZkupLB2oBGFi+9Ct3i0bh5iMtb8ATTY4B3BF0NcZLB8Kuxkw
8Nuar5w4dfVL2kawgyEgD9L6cY/woI+7tCXUDErAEV6Q+xab/Lht00C5DFNKALyp
GaGucPRDcLOlhF/VnZPl77Cxp7rv4EVb1EIUmdbu6pnCX9+gdKmfnZEhDVpHvOHS
ZsFp5eBvIiWMjmBHgL8RCz3CnHsIe16BblgkhZP0IwWkiEDbMeKM7u+ma8ng2Q+t
sLTlcG1jtzH6r2ZSIM2Dp52uw3gGx2znS27bjpOvX8bPWgyHNwijqR4sU8ImLS/Z
vTiAkV0y7CrM21ILTana/+GtwUk08cDahhjcurjEXQS4y9FOIABNg+Czt6JVp0VY
rbkHJ0+JowD94FIrNx3NyRk21BM3reRNJMES9N2zqhVnif8+qfVJXxCeh3BDLHYE
RqR5FRaQ4J4ihU3JQDsJxtxPCWtkQmiQkyqBk5jdVJGcR6R6+WQ8JU6tZI026YyR
W3be6a5Updt6hO+0f4BLItPooRKl5Z1ta1SXmjkAYO+1kUlQHEefL3SmWvx4pQDx
cJ+w4TMlxKPCC7rSrDclnHj3dmlQ4DcEHrdRKljoY5In1NsLUXVR9Mr5ucX/kZyF
80Zh6PvN+WKUh9Wmxhy0u4hy/e83ylLZlPLiMtOVilr+ohlLwMngv6nAq/jB1vBR
sLfHPsHwQqIokG/YWMk/FEo/UXnj0MNty5hgKqyKZXlXH0T0eI0XRwkkBUal+eLi
LceqQ1ElQIabrTJ4pjEnMnu7xxmLb4ZpklHNkz9coKRI/Zf8nHJFGCcto7pMtfo4
spSZPkI5Htxv+Pv9I0afITwA1hJTMJOcz1sbYzxVqkosCn9rTA/AJyrrQ+a/lAoa
ShKxY7aOQwgtS8qvx8Cqo/pmr/IxLiXeUfTCRfTGoOPUn/2Hdr+yvinuB3I8P9sb
OotxXZjSY/GNCylmE7Ccrg18nCm0AOvgV+kB7t5CMGNQg21DU0SdyBQudz3gtKN9
7L48W6yhXRZMCmoGAWWrUDmhb82koOpVVP02l8swhiYXJW/YzrpV6kLAHrsFniPZ
wvQsSlThxDoIwjVynIAwm5ktvsu9LLKM1Syvsa4MtTZeyzyNBMFNBOXHyGRjNWWc
cRwSEzWZU/DA2dY1Q5BP3tWcxdjLatDy8vcfCuOUItmy0RL5U7yt+BE9l6wldTJK
xXPHCAfL0cxGanooEZpTX+M6yOLxsbEFclCSvwnJAUuc71yOoCRGpAABWQ8S5Af+
ADQc+44wxCeF2memvX9lbSdULZHO/4KV+yKOLrNtHP4jmPVxX6z24QahJLPeBW9v
jgkviHAMbtsXDHcSBIUyE841T8VOXdOwJFyzcxF8cXVRjpS8K8+KiBQZrkLNuztc
tn13EJc5dxSne9GWEi6oZPe35wI+CH2ngY9vcUldnoeO/yTzB2MS23ywp97RY4mZ
X3hh9EDDW/NmPYEQj84IqXpbxeAdjUvqMdVJBjVi/RYjcmay1LhPF29Qo/T7L46W
s3kVp3XDr/MWr9GhtOgS6GDNDqaZoz9j2k1PRSv5bAR6TOqdZG873EgZVVnXvXUm
zhgIHznh09B96h3eW+0ZsvjFjr40aifT6LU8jnEsV9lNXCXPPeKB+6r1y5qtWCiY
PGEcmTHgAqyTG8835LgYnWNpmCUp/qsa4pWtwcUUgEky9jBr6SJaMYEnttngj7Vk
VuWa4KkGlllPJS62DI09c30Z819lcaT1yFMf/yQbmJ5+g1wjMM6gkKmTxv6t3CjR
IsuR5V+0afMztz07kIwY7pwcQjbOuE99VrN5AaJPqYFTiRJmgJM9mpYjQpOmcZHm
RNcdi1JgAzgUsFiaCQxzbVFAIRjOm2mVikPw0WVWnVb01UbrUONhxtEDdhaEYmjL
ZgaT+Ryocl72tfT8GMuG7OB5MqAYeyHk8dBeghGgXjwkqh6X5h94031J9J9lyUhm
MQLRnPI2EhAO0XprMilHpNI5BIcl7S9WnOpXhditxxx0PNnrfbgTQUPBEXwVi5TE
FTTXpj8fgaUvD8HqJiBLZa4ZPw5cJ6UoYIVXLUPfmtE/HeZAmCUa4GEFavdqWA03
fpT+jxBXGhiQsT3GkZRS0aM4kSDRVUHhtN9ZuWJTqVnboA9eeEkmg+BwJcaqGf0E
8Xu9gNrnxhrm4OdJaD7TDEc2Ahw2eoIugRxVTF45k7JIHFB2fx+YFyQ1cykaB8sK
+tWy4aCLIo6vko/J1fZl2IxwTD+gNqoLtyq+RO1f75WOiqrPDLczn4bs5BaVnmkb
okWJVYB3ClYJhv514QSdTQfk2OdbJc+unrt/J3UzIDmUiJHuag4J79eBeTnqqdXq
2EfLUkv9G2nMIpMnk2kWM8xWliB96m+vOwjzaGkF1hLfccVb05ARwAhSWmC0yNRv
m6fRr8c5txmyWKHargXIqdL+pg4EYHFhcHpV/PveBSf5VyavGDlHM1vfZOexAu98
7G09O6HjBRS2lVr8XHR6jNF6+MyIACuEkhJZmoz/zGfsk24Q0st4EYCDRRHbYUas
5fDFFG0lAbT2a4sKaK3z96mweIdjwvtbj0VTJUuIC2arzgS4m2NpTzPQK69o2MDq
xGWEdJs69dfJlC6T2MpRHEGxBd9VoFLXewfaBl7kY9ekNwOZ8AXpvi/tYOi5IFyI
vzjya/KWFwk4zg39BJybVvSEnyIscjM8m3qF3l0qwPKhWrk2SMD84MdViHPunui2
cPYZSamShisHr8WHBq1/VEMaJ7JLQpFIYIsJTuDX+Wh9Fp6kY+3h18SLMda4NdKs
Lxub/Ysd1X17djxLUr+hzLli41wfnLlgLxM/2PwtBBxF1oWsNos5uC45rFUE7IFV
NBrmmfN/ZkVSxvaOkRJyGtJuASJEijiqToaTFfmFAIU809tVR2Hox9c2BzF1gq+m
E1Y3z2onyCUTcSqIZ/5ZCqWmZ75R+FuHeleMnUtMNIjTxk6W/TBhh1uM1ozAIlrJ
j36ZrlfJkHUzBHxcOClUmM3Y4FleWbMHBio0mD4suRxnWXEgQutnelziyqACLKzW
L5X3A4od/DBYK7CqpeQruomFTD2I3iugGS8BGyaerZAfJUF0b4q6G4B//PLj5KAo
FcBPYsbXzR2R/qsV+uV0k2yR1Kr2Izz/FlazNKVKOu7scZEgWbq3Y4+EHsB+0O9c
K3WhYgYovxTL3zLLKEFytweU+ke+pB0G430xge3xjxfIN+ak0jIRa3F/415jfFRW
m0F6vWcp5sbwcLf+jEAlGCc32OFjoI5bif7YCzIdk/gT5cAHSWsH8OAGq9pWhoL2
lkO2aTNiMfEqRcG9/XM/fgtbBbKCFw49opwTZSLaayeiacpeclu6aS/u/I8zzbwx
TsjNJ6ou2SJWINh6mvOzqWYkRdTU62XdKAhL22Bj9Ur3lEp87m5UK77Qkntq+6Iz
P0ghC0HiP1Oqiq7Fp7OfZDLl5B6pWzvBm66CJ4dGbozKjqkck1NXhWd0DoO8WcZf
WiABtSZNLhEXAcRwv2oNd5m/hRl9DgmX9Op4+D91xkABuQKMF2EWSBwLGTOjESHV
o/Rbn8GY9Psn1FA/+etqi5SaAmUBNLSRkd2uOcpljVFPEx5Nh2puPgZyzg4RH/pZ
Nq5RskDy/LWcshZEaDJVna12JJyeatJXrcjS5BAD2Xa+rV+mWa19T3vxygVoEYp5
I1MEQAVD8UmytWUyPjLZIKTZWqwSlDMSM6eNfy0KL128R6t3RSiCIoe7k9Hl3IsJ
/XRWB3E/My77NCfG9/ZR0OTlyNruxZDgqjvL9Gv7g8HblVvBQVTWirMe/SPtWk1y
JRFlHO+XZsmVQuDL65ZG3DDnTXLMHLHaajNxifn6aPQ5znLi2hccA83+bU7qotOa
aVdRtNNR/aZVKZ6XKkC+GFjI8Wnz/n3M5G+UbiyBh4dH5SCJG6YPsASGHxVw4ytd
JcQA3cvc7uyV9he+lJjEwSciTZGngMp7uAr0wI8xCgWXg4DnJRlRGvQ5dUBzHCw7
n3tkmWqeOdpiDbFoqCS6OQB+y1FaWpr1Isn2xIfxfxKQgpdWDAK8EzKBSpDjhKmz
dk92Tme/FvWM7pVzK7NqZ1KOllpvLVb9IGWrO3DosP+QeNn+U+debjdOWzrDmuGY
qnM2mco4gyXFg5LtnPojuB6AF0VqLuCRewEfIacJWugNeiGh2eYhOOkdFC3OW1sQ
YqaS8d3Fde3Ge4NZTbQ+9CnUrsQ4dCeLSNzO1R/ZBdowvFJWuvg0jHY+n+Homg65
+g6HU4fVMjvtpn5TQfKKH66HrQEySYiM42F/ws6FiBJbsp/F51ozta55VEWMFwOl
PGu5v6n0dAwvB2y6c3VxRvZufwQ7qRGBysgA2ZeapWtOfaL0ELFjE50LR8oEYANt
6KhkXOyIePRb/1v8xh8jsiEzhXdWWu1QL3yTc5OeuTIiPY550GC3HAbPptJ2Xtf5
W9PKWyDcqD2M/1wUzLBdrgd4Al1eKiE6SzOog5i+5YXHEYh+Bo/NJKZE5RZTrThq
BbFcbOtQ3mz02f1WoQT/8tsLSgyiH23w1vX/keVPjh5+/PzrHvjgobvD1tp9CbJe
hJDY3I+W+i084dMbmcF5tIipRlq530Q2gqye4qFZ4eEr5v4y/hHK9q84CWdHlbKK
ObYWbtHgs8h1GVjs5P5lRunBqzq6NR1vf88n9CtZRU4pL1YZa9NTTasAuZl9QGY9
SJhugoV3RIjk9BV++r7vdRsW61q1wLAUYxJWA/9OX4HK7gSc6GXuUXR6IZT3iG9H
22vTFzG8yogMlT4/j7Nfq3c27HbMcv7O7Xn7ZTnD5TA0Cd3xerqMVu3IsEZAHGTi
RJEsdhNPiHgcPv0G9ID6O2wWHi0I1s7ERsYNI0cIVzxQJajv9EelmAx7oREl0Ut0
pFS6p+xFyb1T43a0p2finBiwN0mtJyYqTBSf5fH/lBcihj0l0S0MyAY1l76v/Me8
OrGgP/vZo26/TjUiOxhjWlA2j5XSqd5gHpWShhP3VDb6wyWR9iZ4uRlWHzJy3/rF
Ej6CX00XJKmDAB0srKFbgd8Kn4hbnZLlOBeHvbn0FpZ29H8LLbGA7U6VN/jdmV8Q
w7y0oB3bhfMTv8IFtz8MmKD8oUaQ6uyYzRsjq0cTWQzTjRquFmZpt2HWo0EEh2rT
LaiI25JDGo5NoCFtB4WFq7oquCe7S7dQqxY/AOJb1TDz8AUcHA5DWc5gL36SIXBJ
`pragma protect end_protected
