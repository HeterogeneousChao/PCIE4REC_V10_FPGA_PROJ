// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:43 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IJNHKz/nRshKI7SXaGTJNn+jqm0hVEa668BpngpGFuHabCa96DWmnaAK0+eZaoSs
803T3si8qNSj9lea0EuLJ9vA8Bd2wVs5d64ECUkaofs6kkubROtfmX+YJlj1O/WL
jm0h7VNpalLHvUqZArXiHFsDsUxpc9JHgTNOCDP1YwY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5296)
d8MC2hQ7QVAQQ+r4MitmrwHi+4O5xgm48I9BuBaCZIpBMcOa1aA6uGdWPiWiM+TC
BOnAFpmB2/eyiufiFr63kKic3uipvagRQ2z63l/Z2ELq/l791L4NAOivqDzMPIGM
Zmcb9C+u+WXJ2qRDsveYP3dJK8Ov7u857nSZHHrhuxfBeOfsCfYCev3NoVBZYAdA
Hhuq4Pd8zPJTyllQU9QyjRr+XMFrErkrWKxQ2+whE7rIwvtspDAQUYM2TsnTlOtP
jHf9Pmt9SxhhwmSUuKSa701+oXvvy7iB1ssOIkqEXanVLnDAT+yJV2KU0kwC9bbj
K+fXfF4rgztkBTfOuJl3lhmxF/UMZVzvSR97b7Kq5qTI62bLjr0CevqIAnR26l1W
ne3UGdSjDyN1siVHP0ExI+NMH0/3MvBJyeW3WyA8gKQa7rfellbrfJigGd03Hy6s
T289vT9ueOHfpva/D33e+53LLEfiuVPJIcdOtU17bYxgcinGUCYGJVdnbkr61ECW
TNfSOnnuDzpZ+BfJ07HSc4nNObGAaKpMmXTdckvaJK+PSZVK8syuhwPeG+TfFFd7
t2CkVnGBox92Qzjc4cricarrsK3w23JLyh8QFJlhM+cFERVhjOvo4HvVlkgk8sj4
CjJprl1jPKFAw/sTZt0J9lI3Dsu5zxZF3gnu/+Ck+2vNS7NKDQx71VPElq+aNgyE
ui6nOn+cu5QCfrb183Mtq4rjOqZ486OnuGMVh4+rMCEIIaxlh752roXPFGdNXc7R
TH2ZzRSD8RJZUAcO9Lc1ilgXGWT0uVWZklt5jgHC1Xtu6wl+DW4Ru3pojbhUxflr
CxqxuQWHTs/zAjuNraHR0lAdBEmr1Xw9/H9Gzh7GzLEwqsnfgy4PAA3Riau4In6m
JodnijBQfwRyvv8A0JTNN0Z00MKZxmIzvNaASBb+lVK1P9zcdrwI2DGPFwsSudMU
WsKRoMDKoUJqn4hMlTUeef3p7Sf7xJiL1ciBODZ9cnwhMJUfRP6D1Jvv86BL4Kth
4fyRvh5MzXVP5YGTeB/WP9CBYkwG4ZaKcFe4p+0yWOi4G1GCRQQyRnR3lJekdIfE
aZLbStbHlA+5LZSm5lYRAO7jD85wtOUBZ3XjIuqh3UCvRiucTgvsblwHomR2FwC9
Pn3466RHyUujY9ISVm3TO4jPyVTNOaFB4ozlXnHH4kbJMaiZk7U8MjevwEpumJiu
/lTH46F6DgW/d1yqOarkMCuPA9243Grn+238hcGm9eIGVuXbSi8QfKpKAiYVEZt3
xh7s4IGOQEu+kqGcChP99Uv/cd5Jo2T+UFZCNQgPCUZTpRqdaEuCvGDdK9hDAl9E
gtWvzNywqE9fWmZ7XtZKUvt+HExX8YbuTDG5jsvTviLCGi+GK7TACWz4ESZtYvEP
JhR1c41qnwfB0Sj2bKBAL4edJHlD8ZXQYyAebtI4grWhRD0igIyzNytT9GlKHreq
kg4GG9wKchQl8iTYz2blOz4Txd5THYpV/aGfVXLPizo/D0WJMe5I9Echv35qySi7
m21XYSVzO2+pYQoiZtmKJpsqx/Ut0/15KFgmlE0dF/lbalfu9bLaydBAB5Nq/uUq
9tCkjfGMoNJ3a7eXvJZeD6VrPY/gzLDZSer8TfAbvKDnbtVJXiZdtgT0Z7e7VytO
Jn5wdfPG4V3eLyg4fBrfRR/qVlOozkaVLLzuAB1zkssn+SboKlJmQh6k7F0yZEWu
n/jn6SAdXi2Rq54NnrzgRckQpMSyY+iOsEK0umQkGV+naTCnBu9wlw7KLx9fVPDw
stg/5X6E1ex7Upu1ir57hrlFPVixg4qBHq6g7Uqj4x5fEjGLBIJzZqw2JsJBXB2E
F+7fKW8N1x+wXtShWittW7a8fvoLlLAg9Jm5eT5HkyNSAmhJZ1Zp1HB5nsqRcche
i+eH87XvOP7t61ShlBQff7PKa13va0NIGJ6wb8qYTWKYn33PfSU9ActBPG6ayBth
2ATzzn52hFF+6OQfQHs+WInBCXtAwL2hj6/+29nenZGTe1RSLgG6Eu9CqpG0cbmh
NE157JQX7AQdlsBMcbHui4lJ69XK9+wBrWSdGFz1km6YQnjNkyRgrtbIxbbqAZS0
bXAGr/0lgwftciy7hn+l/uLElzDSykSveTKuhWRtw1TdHsW1EHpJgyiDhglgFEIu
G7Sd5YtYYGMWSe8wZFy+LSpXapUA911CsN7cAobinu0jw2AYFSCziZgwbyZIneRw
OTyCblHEGG+U8dqT7L+IjA6peXoJqC7zQGoNZfHQOS5dFum0CVvu9WI2r/DaTs5c
Uoc4vxcMj354IrOlcJG82Kiq4GKEcQoXvbVDrcW1JpCBf5f/Dh2RqBUnuZaHPyc3
1qI0O6SGVrpqDypBL0AXCBMnMqh/pDZjF5jOaSqltc/3nU+m3yATFeiNB4b86PeM
i4brb0IkJ7WCF3p9uyV2jvt+QJ1UpIGHvR7rfloFwcvThUUmCPtVbqtZC46CTjWH
B3aAHMtS/Tn85G6EqYNrZIWZEvpUhC4Dthzn4W6nDPLWWItS6J4awdEc/jyFYDb4
fS232W/dZM+4tMAYICz5goKMTZXWbL0LcH++ImpGTZFo1+r3MJkItOSOFIqYtAAw
Yv1v1Rn/ZjHarQUbn10K30LoG0EyBOFysh49tP/oGvm0G2+qe8jorgFCS5/bVtwp
xYtDuYdHg1vzxyBggJH9Z6DjRiuJJYRbJ0oRqHpFEFkIhgbP2EJ/7UMA+sZIDKAc
Nxb1K9pqkhqD37m67LcXMUZokPZfVmR+WrGPq1kbLxgw7rthcXZeKmThLDRF4Qm1
LAKl7+eqlIYCRMJqwa2F8Nwg1Nu7U9k1xVjE56l7Wz0BpHPcJ6IjQIcdqM8XSUEL
eHKZXOBJ2XE3aRz6MkpWtDj2KwCUHw8ki/sHXu0PwxUqIoBLAH4c5icagJjUVaiy
qATEtOLbTChqgMnDOZ1Pkf1EhvVwqWKv3+nVK/dZeTsyvvESuId7LA4XrN1m3fB+
V0txwpqjbhvQ4XgoqvtlOf5bLpaRiDPjSqIxdaft0t1n6Y/r5Ffiw4yt03qmaIOf
5aa8h4Kk0LV0BLQdmf6s3pYjsU/qlPSh49updkWBlCr2JWHX7Ilr2BiXI+rf5m15
y4vOMTmr2VXA+abinU+0JtnA4sGqtGi4BaAdQXrm1Y9C96mRdte3rpQ0ruPQck5a
Xo9/mN/UV7fyaWayfVc0C1vGcPVnj89ap/s5IX8Ky1jgNp9HkB5gESspNp6nwd3J
lIIIvlVTJiD9OV3ifX/eA85J4NqOn9434V9XkbBcPHYl9vheU6wbk4zfHwYGeaiZ
7j2PvuV+9J7zPIGEzrRxkBoo/u5xpFsUcB9nWpfJIGURhlOVDJyjqjLxifJh8fqs
+zm0Ngzj4Pc9pie4TfozzY6ihQxTyX9cUAKU5Abkv38JxMSD+ry2qsjfUWYV/kOE
sW+/C9dxSIUNXdqvFFwCBJ4LrdPdA948wdLKBfC24T1B/TgWtBb3zsoiQHKwv68O
CVfD65fVBGod27wnYJoUos3qQoTq7AAymT4KBNC+z/2XzdyweqEN4fMLGlu0i2JG
ir3y2dxnwzuzYKqK60ySOp8i5Rmo69sXF73lcVWpFkvqH/p/dmRM0PDv3TFuWfYo
RN/N3FNnYzUuSv9IQvtWnYLCPXM7Fj/AgnrGfdSdMw0c8myE207cvmgaV562rZRJ
wtbGR0Z92oSojavaKcDPA2z1w/SW7b57VzYxBKIIbf3NOc4NHslbWgVlMvqwEc/P
ESPSBlvaWRQXBwLovlPcyBCg8qpBuE1kQPA1wR7PSGZlErt2dt1U1UxmSlAGi5SJ
K53pdB88zf1SfNdwMp6dt0IW02C/Hw99AehQH8l94Ox13yB40V913hVDJlZl7Xdq
X7bgW3FAb0JX1jDJ0b7bbgdS5D9qSiMNBFKZ+HKJUwD+6UBYii6Y/y3OClNnPvnE
dzt304lXjhz6ViJPKyLxRc1enVcsQTw/pA/zP3nQrN/8jLZkbtskZErFBGwfdlsc
Za1gxQxGFwmBOcnmeIltH409FPbzzm3/OGiQEuyp5328WEwAr6w6IrUV3ebhpZQK
Sq39opbiNvjK2y7DBq7bNeV255SKBBu2yPFrzA1p7tBtI50dHRuSIja8b9iQ3apa
NsFoiWnrySr67vs9uBRAtF/LR6uQ/dQSNeMMBYH9VohE7fyguKPMHMqG9hydv9pH
Gg/YcDjXPMM+Mb8oSgvFBlBj7FEOc4LnLUpQCZJhKmE220X5w93b63y0h8RRguGu
izMMY2PUR0D4P1CsNwVebK4mjKbdfCRueRpPdkUmhwZqHSN2136MHDHIGrI76hzl
dTL1XIs1ptQN51xM/cv4vYfOHr65Gp6V2MuPp/FCplsrDCTkzTfNgR0AxD+1NoQU
jfcrHX9LLA0HkQoIEefl4BuUbDNlJ0aaH/asp1z2BwmXofadEF+4sj9rWqF7MNOX
i+UzQxjapxu5+h2mpmydaOXS1y286PLzD6VxcQX5gAkOuktvySW93myhzj7UgN9d
yx45lgmWb+IscyezsDliLWQCkARnu1IqsqHh7se4MKuY96Ih9AYxcBk0hRNpO6P4
B94nl1HZefNB+6sFrc+mmo4ZeIbBfMk4+mUAqlbj8AZwZ3iI68qaTUwrRf4TqAs3
B87BiXLSUYmvhli9JRd7SuHFjgLFJq6DcFZDPmDFLj8U06qcBcFXXqUsK3+Rx8V4
WtIHHbszVZQxOy38NhNNJjuyQNxxHOBnDhvz6EPLAu3Hw/pB9p/OPccgpaByqhXg
UuOe6VewnQ7BfmCSKREgaKRrSHavIyHpCq7QdJJ35sb6wrfgkW6v6b/tZkB/oWlV
Cw/tDtK/2GWWrHgT5byAZO8MIIcWQszxyXcULpCKWL75pGpIc8uJyFRrUilcgqEX
Tdj6K65xf/09+3iiPMmfgbD/IZCzky2KfSCRfGgiBX+NOHuAEYigZOQC3WsAuOi4
GuK4d0EqvzyVwKgQsrkEEzdqeivcSOf2uLcofPYeaTrolxutY5drOhhlJf6wpr+E
+8SeG+jkeRsasrDrRu81a09napKk2vUXcTKFUJdVG3cwJq9rsYYxCbgIcirFWqtd
9vceVxmwK/eHsz1AGfNghi9Ya4myZ07fhTw/jnwkiMeeJ0EoRfvaqyiUVUlZB7v1
mQBAFqsxjPM1vJvEiWd44MVlotLJq3Sqlmnu7OnxCiomenZKbZtdP/FVUSi4PAt2
/hAdMruFs0nCOl7XRfd2bhesXg2RDXukjdYHqgcc5aR3U5UDaXI4iNlYEgVnxUdY
893qPe2/SbVE4OMcqQ3/fg7omR8XggRBYPy0gHErgb8OpnU1JUoxOAAv+nX18/If
WXrSM+oMn/eC4HNG564BFSmAMhooVeaOxHPEwSARlZe/14PIAVXKJNuDz7vBPE57
ZS0IXHirNjlTes4jUeVR3rhzTqAyHZrpx1MxQldYMoFNUF9raRDKDq2tvp4HyXv4
AjbfZylaJPkuQHwcUBq9USQtx6+GAMzJ6j0c/y/Zbe+FnjERPH62SWRo7U8l5siO
gxAF/LFx/0/gEKp0Cc2CCFR8z8LmKQevRCUxU3ulMV9loJPGA5yhXIsQlYhWGYRn
WmtAUQtUYfYCV6fTy5YrmtY6rddXcgUVAIea30EkkBbJutconJNMIkbdvbknBA1Q
6Xv1IWqBPOAtOPs/qFW5S5vK4UoCcQbDRGufOGUvdt4Ad4nZQ7fJdGjOdluD+Fzv
o8pmp49JqbOFBh/7Wa1bDMFIneJlGNMDyqwEqE7eSZbnOzW6OR8WLLo7r42Tozko
jzHAYwJATUrrKqtQWDXo0q4OpkhfSQdQ7gddxhaHA81PoqR4XdpLIqE75UGPnmB+
KNzlQ/L5z+XGOzpMwFqMs95X221U/tO44dPm0Fr9IrEBO9gdIrvXu35COx3GgLfq
++fv51Fkprvc3zpZt16yrAV03nMZFWpsvWBWakTMQ2c2c3Tb6mmr02V+6ZGRb/jS
q1Ggu21iTWZzgRllpYYvIF+9D1b5Nqw/vfEgGhviB5zwetKwASrshotZIFjjomki
TlgOrxuzusmV8Sj6ZlAoV6d6K7df4ZTdU5GKingDUCug23DkeZn3pBNWzBExef0I
QgUBDKcc1Ht4vaNHIQ7KtO8ksR3GdJCGpVXrlB9CUPQINGcY6spvxUGSYfY4PMar
Y325Z3jDFxYJxyfrualMkWMGuGvMwufVXIUhhAX7xyPQbS60xfkCBRdPMTaUPcfY
KKQ4gAL4KaRuX3hUF1eEwEkwYUnST6SrGJ7HKx+Bec88BMZj8V8hwRGfNPKUkXai
2McjBOuzRnDc5piDDsgS2OGs8qtnU7P2npO6iXXb5eAHtzvZi5vUT7jVuC3UH7tP
OJw1KzL4GOl1NsHOVCOPoooAhc5TZqGKMWW5wnXSF/0Y7TqYKfArRm7KyWe4AqQw
zg/wy9vOoEEBMsud0OnwgJhqFn1ribJrBWZmAbmzDRe8Otad0B7IHWuZP175nB0H
DcqfmSXMfw21KvakCiQSYzgv23VWYDo1fg7O6F0F0l+7EGSQOAmwLBLpwwDvLlZ4
p7VlB8w3FiGe5oMock8Qe5XoPa55Gm3PmNKdma6Vsdr8eI6y+aWPJbo70AQLpYBP
0Pq4MRcJoYJAOLye9rpbIyo4B+3R7e7cOY06oV6pECkQEKsCj/K9OulSBJBaf4Qj
hL/NbVMGXz4JRk79NJbI47Pd7QPm2sua17MaJ0xhEZmXTmiUMMPUD0OHX/sYSVVk
z7XgI2z8uya8lWwEZOWbUL/jlXVE3GnVwKHjKzWmm46eElNUMUCFy6I9zfN0S+48
xavRO193xnoznPoO+PfTWF+yyP/6GV5dxbObgF/MqMuo868/B26FTHS8H1DBxHCy
rWQPRGD38rKJOlayH0eWekTVJeW5PgkmMvHK52KZ70A/MOQ17lnJog8QPFD5D4Tz
JZbOE1PAty1eqoqfCCT2zOgayxS1nuy3/bSK4AkxwVwMzVvrxmDAVDfbcf7yEXn7
vDN0/1U4J4W4wL8HXyIIsg==
`pragma protect end_protected
