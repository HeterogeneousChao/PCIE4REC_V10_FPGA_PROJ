// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pg5nIKJz4OicWkgNAvTPF1tHxEzvidhjx/ZvfAylDjzAC9TfIAaWEevN+iTZfPZ4
vLyF3aJWqfHpdeyy0FZ9IwoX0qJJ7AX6++F/gmqT1KZjEjIDdMJimVrwjnKR/F74
zgoIoJjsIxi3VExslKc/Jf6jRU3pexST6sCMSLpfd9c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
1NhKz8NAyLdehJlwNyJ0i1YEVoOghVCRVlGFoWtzVedRIGR1Rb3l+Qdc5sSBDgRU
PWrHNNuczMLCN+xj8uZylbBwBQc/ZwK4E5AWqPvwYhg7R1rygeJ/TUcBBC/ZWHfC
g3pGbXMljcpgmuGUPoyz/kC74Q3qSBtotgzGcA6C4Asm7tTtte6zHIJr9OvlwImL
61vuKil/hH/uA86cdob4QOcFiv9ghluAMlQYdsD9dsVSdEeq5pkljdWPp991uYNm
YIvOWIVDwzZEPmBPVe5Cho7ZHVFyRV+l2w/YBrnD6XYEMGc3k13o+qVjj22PXlGd
HUe6X4//jOK0ci8N6/A+P7zgrGm3AgMkydq3iBDd7Pfpws0qmtipyYIFOH2tvxKt
opCbns6QHLEShJKG6p9ECbAKcUCu1ZcKbGtzJ0jn1wjKi8PVK4ZPXYFXT4O2ScPJ
GZ9fhJykL2350E+AfHlmp4LnqAw4ZooUopsVRsHEOk7qpAOxXPDaxLiaGwdiDWoo
v+PiEtduFV90EF0t+1xkIibU8fcmFiEtpvXg2iu2PRmfj2HQqNr/GVRkg2Mw33dB
b7dQtFfAQToKFmdw94dcKC+psN1dfdWIlTn5dPw2zVv1CC+zWcjk9VtZG96xbmCQ
8AWrHOFqYmStPPGBIg83Ec9B99jD0sUbTmmtj5I632HO9ykVOXmom6lhDomad4uY
7lQTzmTLCQmSbOxBDT5kVv+kSvkaGr2LWSgSBlmSWZnqVDkWR48dsfcIillI0f+Z
+KWixkx6Ged48HkIPg63m9s9muUfHqeBH/flJpWmWD7ccILDTFfWmdrlpKM8iy1q
TM0LuJy3DwYFqdInp0hlv1CJgAuCPYWNR9hhSFx6dVvBQBbevO3Vq7l62yLh1gYa
nYrkAzDbo50vABdVeWJcsPItMikKibCI6fplyIwwk9o+gumVfWhToSHSFGVCtII6
5D1TJMOHyI8QOZO31lwrlnAUGfjKIfbOHfSn4Gutx8juczJVl7+0KCdswEEi0p9v
Ff5BaAiAfAgyqEzXxz+/pTUNaPy8BWJ9YSFJt8Xz1n7K6ljrVMRs8JLHNVNeqp8w
CoBtjWBRMMl9Uvt00HcxEXfG8Hhio3fb68xQvTRhEDY7F1NqZYCXDURFwizmSvcZ
qkxLYNwCcBY0nJkGSDgBa6HookIQcRZ3hwdWvymuvwrkL6157OEDRpk3moLzXs/R
64CHZf6aecinNE4vK/4UhELPD6lKo6UGqbgIVuNDzNSGLHOIIywXIlQkOFRLFD9c
//alyh6y7YA0fSyDW/6hQVXaorY+LB0xGfQ7S8KTKqwtn3VZE0x4GHZNe33fMABM
hXfK2MBsllcebwhjJLDR7Bay4gEoRCWJdgb4Jq2wAilNGoa7RvviacneJZ0O/HMw
qR7YFogWGf5SHTumfSwMyuvbMdB+6ofQd7B2Dw/DlfxKSqOL4+DKzFuN6sCJFVek
Su8pjvqEFk3tlcO4Z3P73nSQXXTDkr/3Y6i8CiZaTD1z0oI8QmMQHFEqm8xHEkIO
wqp3xc85xG76dtfx/GD2m/jrX7nxyPfmhfelm1gHhC07WQth9fddGlRoQ/NBMkre
elpnUlMY7nw0ZI6Byr9EubM2pqp6KgmT65nex8KC4N9VQJhOIdbZhpVzbdJXHq4J
45d2yJLvhHLu/4tR8TXiZdGpK82dnTDunFptre6CCYKXp7lsfD0BzJAhjbZnkQNA
hWlK+E/Zuvkk8qSyeB/BS0fyZxEFlfTqkRl7guW7NCaH7T+1HdFCMO9k+ZMpQy+H
BRaa5fn1bLjCH7gyhD2k5sjaSzc5Ix8lqCUCZM+qpeMwgMJwVjXA9e9jIRIFgsFQ
UjsBNyM4EBAYi/2ZpAzqMrwn5WoJYrE/yN4PIgd83K4fn9xedFveHr4njP5ZnjTE
jn2ai7aDpvYVk/Lh7c/mJpnAV2VuI8HwBZMe0kw15jkratJRuE+LudAfwZkR4L7+
0mDHuY9U1+pF25Dm5WZD/cVKlvzHXF7dxSGnqPkxkinhodGy4QTfywSnTywfbgAL
Exz4Q47ABTH4Bi936ZIo0TgKdSgfNRB+leQTpXzXf7IPpXe+SRKkrPxdEwDeEyUL
2qRqdcE/EF8Y6SkW1ZcSHvlCY0kGGs0YrlVXV9PLMmDajlT1J3y1912GPCX0eum5
1XRShzIzbGjKDwvh5fDv52tdxdD24qqMKXAUzwvV5z9jsedabWCMVWJH+ruue9TZ
ODu5LBXb4BD+XGKeh3B07uI0x+3+Ff/+RyWmw7vczzZEZhDVS65iltmX2i9KMFbQ
A9xHcDTiI4qkjhyAO7ClYRo89KyAuRzcL2dvmT9CUbXN8cpne3zNiwPto9U400qt
9rZjCTWgdzrkPn/FFOydU2BLB79o3ZTzvFJBKkgwYWrurGD+4+/Lx/ttV1y380pb
an+YUIOPaLoehGiX7uHSLSPrcvW4NXfjGBLqW8acgpsgH645mkwvqboyIgOMhkOU
YTDt6FDpByG3CHoVM0Ods97BlG7NRQS+D4Y2/mzlccwNmRYUSd/DVcc0LRYxo29g
+hZePu+LI/ij9KDa3bN3DNUtp6JtIdBJlCDLwETmsVoCS7ZWpvfDUnKy2pbxJluU
dU8ltUTgsP94uwWGTZtrohBj04rUtapHti6p+1VAimUwa+flZsN1Pa30I6oO+bc+
NpQGEkEtTq3Apg+s0iqRM2vK0ezydMGW0NTD3BFc0QoKBAxj6i1q2IUAL2mAHDqn
b8axaJJjEGft9FB2KIb7Ae4H0WJMV7bxUHXmFv+IxL/+PUk3HlGVanxLWaf4HZ0X
8fNFsIrNl+kYuIqL68EGaqEmm5NZjssWWa5ubQTxKjDi83kDHsO1pZ8EKunYKIdl
7mAl3ub9oJWcx22quOtPlQz8hYR49+/5BrSZ4bS63JPb/+scwJKJmymkLbthA6H0
cVoGsHkgw4bsYkNyOM9nDdSJp+1sGkrn8gTRN3APrksV5POPO5pJXQAaMZ9kxX8O
YMv1S+AdRXm46spH8iCcdos0/nw3TgHKJZ8CjW1bTDLjryn6n3BFp7vVnKpM5so0
MhEbVBGmEHQTnTixynCKod1pwJOaxz544Caexz0M3AQ1FCoRBiZxghVSilySZtAx
g18A61vEYv9U8nV2utLNH3x++TALdpmrf4JNyXDkJWXOVUAZkEj4YPT3eMeV5wo2
BRhXXq+EjvrpqVaORR/m4rSxuLm6hLyrvElRuWDyh4KVVk+E6TN/xvESt7wDoFof
bFtEaMuhz4OKEV33pglphqHfFCMCeORREHpP1tDeFcFn/MtzwxQnKMRvs3znc48N
cex/dN4KoiKhcyZ8X2aCaSFd9xcqSm9eAXnP2KCDrdqjzp1PjBHfYu7w3ko4If1B
pN4L0V6kJGt1S5V1wkvxg+d/+PyosESpdKBfrqkGgQonblC1LpDywa0rb2ZhugFy
I7yK3VOkQba8NqdZIKVqDS8j+KrpKqSE4qIOJUVoxmAaikoHSCVlllkkXv4PM/HP
QxR5g8CFSQG4vfBnd+xtrSqPhV+7/jKUGdfmcF+69IvA4SL+5H2OvWPiq/7WORX9
o8mNUDz/1xNshJMtA/tfl6NfYe42lYtj0Imr16xSzFd7R+o0YydWUpmutEbReitA
JD9vKn42O4UQ9Ij3NqizA9gMz1xR5rTtKlYN4I9X1N+mmHTMu5eCPOCwlhf4+h/l
wOCa63C79oGA3RAG9Df0HvnizBFWvnueLU6gaDqsy8E1vBXX4VVasGUbU3c/0Kay
YQG+/eK9UcNfw3c65MOxLRlsicI0piiyHs886BwKTky0TwjBCHJMr+CX3SaAwyyk
wKK4iA2ZIxcjaW1BhMp/oRuXONYDlUiD5/ctNc2Ptef9TF2WoIkWvGktVA4LiqEn
ToOPxVthADz/ZCJtFynoAYkM+FxrMKeZT2L0nxmRrBgEekKP52iCr1KloW/bWuBI
s4zvWwN8RfjEGldiQHVDJs6TxHykZajCxQYMw6PUnESH8I6+ELHIZD9TDRyYJxKF
A3XErXvG8RNPvorTdAcgCDBO1I1ZZiPkbL/DVNAc/OQ=
`pragma protect end_protected
