// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:28 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PxOqScmFPPIKK0Ot87oOFkXv/E0gb+d5n46nZsWouY4V9anCC7tYzZugU8n5Vpx3
1e/viJHKyNjMMneVHe6m/2Zi2rrwpX8Llf7v/x0CkZZ4nd0fJgCDY+0GFVs/OipY
dUybpcQZ3Vms0Rz4q0HcVGeXlmcNtDGRmabyIUi0kM0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
zWG0qs3Nof7ldJEOdMarRx61qZ9NCcCD3A9ulOP9azHQrDlv+j++bRgT/wFWxwFl
8NTWMZgmpX38cNfORpvdpGetx+wlQDiPDZUx2Znt4nRE6z/etj8+DgNjse89jzB8
LePqa7d95kVkMBOEvRPG55c3nO7G+2jKKEZtL5PjlNVGzKHCYR5AjrDmIRohNLmp
2mXLInwHIfAz+5AIo2MRIkw5vnU7Q/vTrmx9hlVlC+zgP585wpVboEd9mQ2ZrSNq
jmoiI4jrsTeHbpaJUTuPmmMFjk/miJTib7pIBEPAzWQgoEatRFi97LEjZgPggqXa
iU1TnQm1bFOcK8cPELePVWXupZxwiFyvuygVtZvx9cF6hngueo33BnLhhX/3LAwn
pGi/P/b48Uo6MX0fR/e73JcB1GkC9mdIsBN4u0tN38Q4jqFjkXT79DeUDH2uMa9C
1zJqHUX0JN8dIZlDAi5s48/PqUg8Gt6VM3YkdsSNiBaYhVCWdxvqdoRN5HZiDDYG
URRtJNTWCA67q0l5a9jU2zWhFaETftVEjUepL7fdGwybNffCC7tRvfCTiyiMXnds
5bFGpM8tLuUVLxWxnKih7tuaWuNi+E/5aoDb9ovxQh1Bj3pMKzlYOKp+jJGTn2Xh
hMFN9ad7yAA0iGf4bBO8IZT77pZ5qJ2Ek2Xm46SmKNfmEoyEgyjJogK8kAkX+GTb
FR8FQB4z+gnc1YZ10iKeo0WdLwWtvnqQXSrRzAIxOCyOG6fdcgg38EkG/6HN1B3e
vs2h5Y4tIppuRbbqji2UKYMIBXQREpmObTPATgzxWJ49gK61/RvYMoAReW/TDYrq
09Pa8mGNeto65oX84dNgk176kId5F35BDhBNvWlHOgN93/BGDp6PIgn1A+o6G7nS
LcsPAhLl9sOsbqgPy7zcZryd9YMz7WgUSvVCDCePVrQHTN664tK3Ra+MLQ5MyqU7
zgx1McxFcnlsDZ/w2qf+qAILUYhYR+EuQAC6u6YdQTENeWLYCaR8Oocw3h6NEVgT
lAZPfdJGLJO6uQgneTh9x+POGySN/RcqRKco++UBC8UMaR8xbS9Cq+57A23i9txN
WI5ff/+MsfWIpjJLvIp6T0jdM84CwxLUlbTG7NLkvFignRk6gL8cEoHayJRIXFQe
5w6uryoVIw5CTZezAJSbeZB/G8JIMMaCHSUjfb8H21aUhWvHawG8YZCyQCdLPiR3
dL39BoQT6/Z0vpHU9X7wbroqQMIlnO2EL05VdweA0wpMCnRbQKKGj6aFabWpWBhm
cvMYYOfsnmA/rIfi8v0QLmcx2G4ldGdjgnr8pg3IzWssdKnRuQloYpPqibwhYv7m
OH4ncNBwl1nJhoLZyTshfcjmVUanDHj07EeSp+Q6qMY+ahXlyBi6WaMLlct3ZRlI
+Dnm4MaMA4O6aWM/7+50lz5CxGoZU3gUtyMoVT/8agJJjBAj6OuZLPLUfJYmRjHk
IgzQSDaFaDWP0k/gm6q+NkYylYlBDDY/LKLkY8V2GjqnFpohnQyAg1taDbILmGFY
MneJmmBHtO6BxEKspaw4/whSH6UkSofBRtr8UWP3TPTGtj3WjvszUobsv9zn+bjg
J6o0tR0QzU3SDOZuhoaTdVi3R5hWurYa/KbIckYCEsJWjYq0Xry1+U+uDzJ00BR8
sn2amgBpJL84hotTo+l3IzM6AvidaKPcSvZbzH/L0LOCyxFYS+eZdMgv9tyYo+QF
Gnri4FjsGzQAbQ2ZxyxsTd+H2xcMCxDgLkZ76K9xa1sqgEFf8kpSHExsSCyt0coN
j9E1wJL5YQx1s+eJbS8FQ/t8Wpi+ZudcJu7yuGFz3AXtnuB16UKDzpl6PjL1LdTt
amDZdkwBIejaqdhhGIKvSbOVUMASx+weBTkRXZsS8ERO9iZ/8kW4XIdr4/6qmDS7
cDe44tP2fMYmn6TucpxRPUVBtbQadDpTHuKfF6RZRXRV+Xblx9buvwNGAEI5PYjG
nhUo5VH91E3nPrRx26wV/kYR4i1OKA6RoLq5dFTMqyae+D2txlCpHB1RZDc32Uhs
I26E/cShjk+JgKz0l5ogexCQfLWSZ56SCFEIvaAUS/Dn1L0kOeF8E8sm4ZHuWpTY
kBZg/2SbuoM0i72pNNhl+nLQwLQBG6FdlmDkh9PvR2Yd+qmQ+LM05iYKx+v89vyD
FMvWQw8/eOBELtr2KEn3r5nuncJCivG1cJBxBDcungx0U2gTZbJIMDMUuL4bQTBo
NyNeEBTh3yM2qirHcISZKKpLlkoQcbTvm4tZBAAL5WTxoF+PgZ6dnPN8mcRwmmwE
0URxuICuGES5024mKdbYl0bNVTmCXGwLvkcMxp5XD0qIDD05M1KxpqWjLfA+IZaL
nHeore3IAqHKzinxkPTXBOk+kVw/a2RAsyrNlPtzHx5cYTDuNoOfs0CxyfihEfau
RHUFEuHa1rcfwPPPXkU/6xBUDdNhV7MvNZNj2k+96NZLD2DFYqx+x7e3JP5Hcqf7
yY3swcdPUnJ8wpdM1Dz4J1vzCDNmUfBDxUYil8tAcJ3MUck0ot/TJjJsRY3WValn
uZHKt1YF3DJET04+EeP7X88usieX0eVWZD/UBwbF55iFdZL81EBT9H5dOAqPKZmG
ZA6W1uvQmAdrl2U9jEWBa08Tq38EY94ml7Bn0HVIv/Lkd8mB129ZKvX5qvPV1DqL
0swruv2yXXcqnjEOf7r3UIRyXz4RZVF+RswI4PYs+wvqQ031qr0KpP+po5o6OtEo
/odT8X+9qVIe86+Gvq8kNpgiQ8Sn3z4iAQYt4/t+VE3eA9YHmWzVKya7M1egkH3b
xvSnovRQLYu6c0KdIagqLL8n2rtaAKz/q4Bn/ZLAqKfkw3ZQrwgbDixPo4/DXVOy
S7luJr+lWhZdGMpO11jpHPfJ1YFXeyeuujHM7aYLJSPbDk7lvE40JEuUU0G3hX7U
QqodsQwWfK/LHsRPXY273qVE+17pWBtxMiSKiXzRqPrNNhLmGVx0SWXyrpzTpyzw
koSFXkO4ihxwRHSZ4Hdy7oTcEcR2eBzfVwGp3fuzSTfjxxEuXEGAYiKwaRaxMTic
oZF4JUquEFwvGRqG9zVjvPOps0WECZVId54ordCQo5hd4FGDEc2dp60qWVYFFPEU
gm+3uVSNYgiYehX6SgRoyP23i/DBOSnHqc+0CftHuY3GZ8sBSxn5iRo9cMzn4PA0
M1LEbgN4I1EdwvsTIbj5G2abUD+dKxU+pRRZzEGWUYqshDYhiKN54tJANiLIEqUQ
+f34rBvwJrhmnyt1bVrLHVv5RGmxqwX+uOGNx+Ft/0FlXQAGN1CS/hK4OxLSl2qm
7wc8EU4TC6Wn9p7MsmOCAl2eSDdY7fRE3QqQ+SbUJIy6lhBTsoY8BbpHDQdPcet/
2TqVHpFXQeowDCM0GmVzC5lvlnWET/vNUoHnHmSrtPUWNHZLR5ddWGnsoKkPffJR
/SC1eVRQ6L3KtDjaWrKxR6OeIglP+hAjo9E5ry2DTEAIilU4mbSXKRqZhRHruhHf
AFdtEYPcY6+YWbpyN7IDX83VMkPVO7jh8BUeaeRqOt5neIRqQTeRAwgh1CsL87BD
b6lpugW8LaNNDxiao0IpBaISL2CaAujHJbpdlHLaxufLO7yZLWWOozFnL1hU6ukT
z2IENngFhF6EllKxkh8qqa04zmvgCnRAn4nxBIoIoxOa0wT1IaIIF0rZEEZye5j+
8QbOln+zxvA3TikPzGFPATFOwdCNkKKiGYsPgw68peFanjWF1V7q2LRPA/pcfj/n
ydC8mC+7xJxcudxhZh3CNw/zs+hnF6i9ltXGN5GUv0F9OImUEzBErz5aaiDOD0Lk
XjRk7jbuBiK3FglIG9EaVvFP6GkAC5Jl1kKK/CZoFLFol9AA3RYadbjGEfazs+fH
QYRyUv127+BlWVMcJznoFbtj3udu8Au5pIgLHd0HjIlIczi0dZYn5xElidadj62Q
46ViOx1MKoc3MspWczmbq9Z+JOFx2xCeSrx1r/Mi/QgAk3o9T4uwRzAux2jGi/U2
zhiZgbfMvKZwWBUIMc8MNOSSIRPOkg+d8VClbpN0niZIZurEZPBnD06GMJGJa1C+
hkb2MFX44W9I31jO6T9OFHaMgbELYkOHHkeQW9oDReBxeJ85TbuR/thiE0E2ipSh
X3CS4a6IWGUb90GWxMYeYsYxr6yFcVati+H/PGgQ4An+sKrTLfFNyv8elF5geQaV
4BGSzu5HFmYzp26El3Hcb/oMXMUXFcE3NEYoq7T5bfp/SIgRhwipPQ6Pv/QJkXvu
s415Z2zYLKmZhPbO3TClPmEwwg0LU42UozTxz4SiRZMW+Qy0rQuwBg+OPHfkPpTj
gC5u8rmfr3sZoSdQ0MAfSvIjBZKLr4v476sM24ZTY2yiIhUo5QVRbQYPkeTpo3ZU
PnxWRbyI9KTQlJRr5x3PAv6Jufsn5xsHy0dRo6ZVnzHnGSMSN44WGwelvdp1gWGU
aooE60gSWScCeQluE0HI8FrzmeWFdalJ1Vt8cKRGc+6f9wuMnLDyJGPcoIPJbqCn
fhYMtX9+z2YuWkEhReKmLBgo2Y08jRvIMy8rj9Z1xigKgluseCKij6WbJ83boflu
HSL+a/+LqqOQUNUkbJnPyuAp/3xawgTeGBulHOKkT7GWz/SN+oCrJ3SFpmswgA05
Avy1zdKqDg5ebA4aJHyh+0OgnhRw6w/lu1VaGVd+cwS8SSCIUY+/dgfMvvycKDHF
iS9cEZ4CfwqYq0DetSfi64XAtYS7j6Rd2xAC4XqA7QoCIyq0CFiQFoi+/aO8rpkp
bpt83pVIIw/8bwiND+tIIeIW3TC2hG++zFU06DEXHwv9oc37e070t+dV1cm2OwAz
+9dKEUV1E/YHe7rNFfzhq5yJy5zFkaNa+LoT2/hpxveNJspp6hF+gYPzDDGUoM1R
5tfQQL/+WqsMFszxUDBIWDAiVB6Ai+SbubozIvDy2HwZpHHdJOtCDZhtgjoDkuw3
eQA2lz7EhR1jKb49NgKSZk4JmrxSXDJirU+xHRvuwQCw2sbPeTiWmq24Ov6Ogs7N
lZPbFJnZPzlG+UlvxqHKqigURjPziQ8gs+hVlMmVf9dnfcIwqHb0LuGCJ9+XDtCa
BgIhiQbG3K56DUVW6H92YrJYZfIIiGTJzpE4Z2njifpjKkKG9N9K5uYj4uXLHs8t
oqi1T17SLlMk+vx0GxmzwVtcsp0IyguMoONCpUbxLsy2n9lUT/Rvw9qy/Iq7pw5a
qznbcCdeAgXRj8kOvcQ0VCo0/fuLtCr1ly427jSxLmCmBNS8drRxagN4Q/3hIQn7
SAsK9EO0QXQElWtD9dU9MykVg74ss5+oB3TksoeI+Z5H4RcqQtM39glQtw1q4iit
gSODJikJL9QTs2j1gGusk4GTfk0Hwr+uAi/a8D/Nc3oc2eMF6gDW3hk1E0fAF2HF
VxH4kM+UFEFV5NfYK0BqvK5OsILXctRtV++jdErVusj7XqpPKCkJByIBhzMBF1Ft
oEgyRcbzNe1dNm6GmSDfSLMGPZKToZsOX++cXOaqm3iADmbIEenWm2gw2YwGkbjt
iCCiDp0sHEux0x7aKFwg2tcBx/oZaG9B6UqballfE85Xx0gfogafkRLVJMRYCNdQ
BPC4zDL9EgnbqsoS3Ws7eC2Q4M/tofHdICzkSnhNRSGbTVZIV/YF6qUN9OQBvk6a
Zc1Ru5kkEt46wJ7bwYRgw8q53B6F5D1jW8eqisruqb8YSuOsbaCgjdGKEYoSMY3Y
2a0DMy+OIABZ1YbRs8sMtVE33bR8OuoOBQ/b2y+770wGX4a2NcFqmLUCk9IvfphV
fRUg2sWy8G8xHZSzlkA08cxIoY2hG2IYhufOMTDpQZHnFuujzh92k5u6UBQsPyqv
Sf1ZszuDZ23Gul7dzVs5BkqKhpsArgU8pOX5RgtmbZcEA0byhT0voE3jVJEdura0
W8nROyJrQ2pW2UGNVRrUwJ/lqriQYtMcvHEhBCzCaqSYaoyzTiDZqf8nkwFDFA68
iY0WuBt7wK+IylQnf9txXWkbrzTTv8QJ1Vv7hSv0mW+Z2eF8/piKZESmjqNHYQSg
eFzOTGAnXYDuDpEkd3AxDBUv6jbllY16ImTeBzkOZZu1fdpZrNC2XUCUZvU0msRV
88to91IxGUA2nQvT4SJFbD+GhPlTTDq8HJSDIopxm3vyGpc29FW+DoWME4+DfoWL
ZArjVphTpz+3jRA/tqWjakNkxGNlMPz8H0nLqpZckd0bj8d/0OI4RKhF9akZ3qO7
vZJGNqmq8Dn4gqtyqLhAFJ0LskgEgFvJU87cDNhTfcNxha1TheM85EMN+GAGl/yD
kQOjWrYAunxx8PkRsocpWgwLL3E2WYMGrjddrFmFst08h3j3wsrNt1kUMD8T7rnT
vqS8iKtjAkAXmOWWtvlfaSnr4IaIw8o6GNSEIskJyBTD/WNmREXPqEINKEz3vf3f
vyxLJWVG5q6zSqpf4iyUYJivofbnxidknGUpVOHEpm89ZGlRb+7HvPeSupVQ1zEv
0pSrz6lBbe3Ib2LFz7ac51kF/9pHDjbL6+V/RLpU5Lr23lyRf7fihm9S59ECwIBq
swr/X2r0f4sjBuY8fI8obggA1ldM9tu6t4xxjahyitv4TJ7QKcghRryHOOMcaANX
L8Pb2Xjolkb/BHCcow8I8510iPxPYDBxKHBNdVWv4nFiUbODezK25Vi72Pu/NNGc
DyRI5bPPrM8nTmyCVTrUfsMXucBFy3NfxdZ0S8e3uyhQFyibFwsarqzfxD/mC+vF
c/or3A3Pb8G4x28cLfnjSTgWG30q3RPhFS8ltOkyND5fHw0YLsGNXfeFNgjNaYj5
c3f5rAEpEHqMBj6zz0MW2v9YqYWPB8chhIY9+xglf1x+CBVk3M65r02L2x6gl/GY
gYmtFqiHnvC36iAxktquTeA/61o9P9LcD+48Oa5jGtytm7V3G+2tNYWYPTqLMqIQ
S1CQoMjpz2v0CM9uQTfzLeiAjIME5O4+CXUWyVxUjT/O6B0j6xUjeVZt9dMLZkE0
o/s1vr4Rp/oJYeBD6S1Ob/29GLIFMHymknWfztJvXTjeKiUKhhpMQguEgnAc7o0n
dNluk0TmG7RYRDNjSRSaYblNTz2gBzYBTq1pTODq2aet50LofqekWUPWbufIKoPe
noC62CSl70sGQ+4tgFyz7TL+A5d5zgjFwEp0A4dGWuUGTEvo8MAFZxPVeiXp7ePX
GG9rRRDPXiG7UZk074nMtUj072Iu5f89bnMekz/SJ22kQCdpy4ilvQOE3EpS72vt
G1oVBSNRG4pI5ejyhTinBaiAeE9BFcP1wYkAb+J6fcv7Qul3JVs8OXe9sCaMNeLT
ny5Y98m1RGBfh2jw5B1ue/xbxJm9czwtoQg9sJ4qFt24nAW7hixRmGgOmMBA8BrG
wTrvlf7cUT/W2Zu/kCBI1iBRpsN8n6bqd3qLBMZKb2O4dTSr9GrEyvwoBOr0qqdG
qgptsH2g8E0gFcUq1LzcbktCnVPDsSxckubkBlC1Iqtku18apv9aRck0RMhywlZH
VxyhlGd50YD6t2Dd7BtbCRyhutvx9Plx2FLv4cwglsHBrW36pZy7wSh5NEWozzZS
0Vp7MCodG4rTl0VqDSZuq+p5KovkOe+Q0yCTMoIuZt+4BOC1FkUN8BXWXVRVLik6
l2TSnyFsB1TxBrXuFYJEuh1KMmymYJe9iMqYwOJI5SS9toYWQjmOruOTEjOI3HRI
spMcxdAOnnKCSSrzJNvUFp6LukUxrfmlq+3jzq5ry9h8aGwCe9FyQUVEriwIjO/U
nstVq+RH/0yBZdzsul5pQooExsiE9R9MyWd71zUHV1HJsEDsKARw7+LHuelX+5r/
jhLTgNzUFIJBxuaUiXIPaJUChkFW5FwzwyAtjRmLinR1ZTwyEgLM4eGEdYaqfIa3
4bb2MdY733cQ4mqyUr7pW8Ku/74pEUaL0bWnFPNt0rh97nL5oEXaGjAE2FDJI42q
OTv2SP7eXsqKPCBlwKNHBXhMMFcQVp8xDnsvAyrigDUoeOC//VdkE+6KU9XY7XAA
y2dCXLIxydF1pa1Wi1Sl51htPIZUefOBXKVAs2JWDvYg1uTX0MH/0mJYhde+/tTR
t5bxcGiRCchnoIkjs/MiqMLN09dHSOQdbW8C8o7AzFwpYv36tY6ET9vx4tLRo25X
Nlm2SvoKLvpbIeVNl3IH+wplEbieUX+JvEE/dr5cA22KH6nMKp6Ooq5Aio4JtIZc
XgFVtm8xlodgGqeu24eUg9M6LBG28+m/q8RI05XqDeACac1v351rq3LJQPe4WGJN
Lxjo1t3Tq/HI4DBJR/baR+cmF/4e9pUrQ0BTS56aekMmRM9RdAEawoeWSnmKmwEW
ujnCcAHUmhxjxyirI29DNE5yY9bgAe6xn0BlpEDPaROtIqr54ohF9N/LakzZoqz1
XhskGBlptE6CANgTmCpFHVtl1ZFD1jr4zgWz8s7oVnN/6P7wsslGjsYQypHtx6YK
pcNdbx2ZQhZ2JrRpDiJgmjdAdsvZrpDa5QR5QYxTBk2pW+lmfwgM/EIDzcQbouBh
XAdiglkA9l22nkvAQ7ZAhqGvLp4kjwyvPyx+3k8EqHWJbrg3BzYskjfzRcyWFQUs
IbZc3nguR8eCoNx56SfEo+b3Hp5hDLmCDJyVuRR1X31DlBwDARizqUl9KUTwJUgW
tYiYlsmmdJK49KOGoOsFWl0enPmRdCftDVuk8Y0nWn82dJSboP/9uUbccGysMCNU
ONdIDauthLKCZX+F4W4xEY5rSavM+hdclZMCptLacZsviH7LRW7ml/jEkhzyy435
ioVL+BO9pnq5zBXC+v7W0n9If5JoL5kc+HrJ/WoF7oo5gtb2qppSbJf2yFJ4nzWt
1Fr2Je2bZIbYUvgoXzFlFAJtqX1TF+Y1r40tDyFESvAktN/3aogHG3FKMDp8dM5H
+xxL4g6Npbr7Iq5morhAfx2Wvl46OuJsf2t71AoxLxhZXRyHOOsq5Yd8n0AykK9m
wzHCIDvegs2khbsj9rtdsoszR7jb4Y0VExynxD3MgeC/BhbVbBwqR+H8vVlcrfit
HAZwgWA/ilJe0OJwzZUSucRsvMqs4NQ159bp0Y/M4xqmJmmlwalLxGbfWhM0Hb/o
+Yttq75NGslsUOv02GK12H+H+U2DrjDSbY54fcQ0tD5PZD7O9k6s5yskpvJ1VUVP
ZIVG+2psrXELzb+uWgsOlV8cMCI2DVSCDlynfHmWFD81CPcYSRQY+A4Pzdb4gn9W
pQJvdy9enSFTdZwLaCRahdzmTX0dbJktLC2IEitW0kySxMaGJ+7G9f4uAXwK2Pdj
k+kNHQPY6p4D5BOikuwwtzAOSsRZFkIFanp1F5++XU8Warv/v0fTZIq04ksCjTRc
+bZ+69mKyKqVG4bWoXoqKQxng7Q+eyNtEI3IzQ7K3+2vLx/0aZromiJmdulA84BP
hV21XHWt31sFPvscrIGMDxKXn1gr/eSP2SvHKpOR+BNYxoKMwtNyGeffNNPCi+A5
SeL8YrqsSeby7yJ1s+1Tmy/dWk0kDyGn8MGl+HWTZlXQyT49JQ6SBnX8h/Pjvfuo
mGJuKMvkYdBu6p7r/qcxrTDm3KcwKq6ZeH2PDedLO4Zh8MwzZSuV30AEZ64DJwD2
0TxRwUivxxTMsFhV9JKBqP+Vog2l97F8mfQT5IfNLsNo/zuOOxyXCNUKKVS8FAda
u+V0KKi6J+XHrfc/awWUBo8MKEC9gI38nbcP6fafGmzYvszgbpd/KAPsHAe5l655
QD9IVZ6lkOAg5LjfETcbhl1DvJkTuRau96VVsj97LOYX7pdmf9TvxEDBDWVKw2BZ
JWTnArYkFeyUbQXmhIMSSC8DD8GBxQYmcHKfEBASVkWO3zsw6ADbz15kBwQ/wTQP
iYb4Id3M+4E5K/N2mWb0fnmRp0wPmNeHnOvUhN6EBzuCgvPhGxZ1ROolQBcm78Zw
4cx9skoW1iB/+EWsPAmZ99Z5oTAh6ei0bqTADKctOUDnYK8lhQib81N8AdnuKx42
AevvpozoKhq5JZOZhElYlz705SdEL6UsVnEe2sbd2sJ2wQA7UoNfOWZBcXegIHZ+
KBcS4W9p0z31v3EC8Exr3UgOf3+IUl1UfqHOWcucLp5envmaKM1tga+UX/RuMPEo
xZxpQI8QbVWKt5yyMocU3pfN5buLx9MmoFAyLIah1XhrKolznwW6m2ttOTeLYMfT
zVXG9kvN6lQCpf0bonW+THRC2OX5PwvIQ13+My+bh34PBUjMQonxLvjbhS8Cz2ef
qNgXwoiCzFlM4FTxcG74hSgO1Ki2ZdbWpC/DDnd/wJmxzlinFuz0gV/Nwg08IbUc
UxC01VfIEWYqUnh0b6a4YGO8MvWteMfFHWbNv3hIRiOFKoReeO9ENkM4nmcNll1F
Dv4Wt1UHTcIISu7/U6D2yz7lBw56KocbTY5xbNewBsNYvTwM9u7zQD0SCj+rsbrG
ga5JkIJDsrBy3s+9+g7diBZIejf/MOCkgq6j+rOwuYwSes/zsTWbA7i9dctP/EO7
QbhLmX/eZxOXc4Etx7BBq0Snp50O7PrQKTg6TcX0+pGrDq1kt6Nnb/40i/YKO6BL
AmOi5RDKw+kIHza+6fO6RHmw0YeiuPnNVuwjSCrtUqdS4TK0A0ArNxJ141RmBVNp
pOuj4kxoLsEB2HyNT2tlxqF8gQ/bxot0QOu/sdJqeYnTWWEcq15HYKTW+TvRv/KS
02a856P3bljdV5TkH4qMjLwGAafExV/43Aiyz8muLUE3YSrT7qjncvT7UH5I4ENG
RB/SV/QXQHJYDM6zhXZ95dYAAo/RS6uVKp3EctQFb5PppvCPaM7HiV36sOhn4etc
NUVCz9d17Ur93FJgnTxbQIlrLuG3B456eV1unxS0sX4cRj5NJ/+SEdbWloiaj21q
iq9h42fYpNMepU7nDAYDqkFRBxtVy58eqkFpzIgX2BPjChdCTqskJwLyigc5kc6R
OhJzWggncrBhj7UBTdDvaUINqeGkfREpCxNqmEsfXvmuNcHP1itO3bpUgkfn038U
ydkKueKnTGa0bU5j5/d1X25yztcpCBV9xW8VBCDuTascBdV7fyOu3yA+SneZrqiP
8//4iOr6MSvxV6mSTCYMENluTBPANQpxjXIIJje44d0R9iN+YznLvJ+tVZE5YShY
H+NQZFx7K8FY5ACeCmyMdgOnhyOx5BGADXeEB7yhsQpHK5lLBcC+4XI1Cif7dToM
BYIug9fKJD24myB8zC8iho775EolXJsIFfKq1n+vJkJrcz90VE/Wf9iKw/na+e/k
wmhLad2R214z9EYpNLJCqTlCmR69pjsUkxjQHas7HBHr7aqRThjqPmbHtvw9TKXb
2kjIUaagi1413kFlc+RFI7tMASCV5uRO6v0q6pkSS6r8Xc8Q5JE/qkAcnh8O9ZQP
tZgp973p32Ko8Lc8x0F58qwPgz1eWL9SHrsMNQkjSrPNC9kSC1IHfFFrNXyutabB
1miPMoERywN0H1p03+q47ddcaw78thwQOQTmJqhi4aiFQZhMbWG93IlGmcbyzqCg
AC34AUN3h92H2xVsj7ryTgqOJVINJISoeWbyUf3F++M23oDwQfMLP31RYGvsMA3c
1ixXCf3awg4u2ujXZJmJbjz5LgyA2UXz0xqD7IXpgOCPzoZWXqV7fbbbTaixkaVX
+5VeshxYByJfMVP2YBDwodlw+QQarMo8BlWfxVTqn/DLyKsojizWekTokvdoAe3p
FNdNmGEVIDhi5bFuavKfxHBr56TIXH2KA0622K/5TpqoFxqHUx1sxfMqjQWe8hcH
afGVWBd5Slglcyx2fmbEdpaWSBqSwqzY3vfe8wovUkPsoiN++lpQKA3b3w0KIq8N
yIydFLUI1RQrqJnCiDTvbvbnOpHO8QCalDQReuMJrmnZf+94EW2kQaEqCX9Uoymm
UAtqmCWOY4SAAaL8Dz4MENdHrJo5a8k+uFsYZZws1eA23zxNogUxjzDcEyRqu9ka
3PZa9xwpwcHrhiJai74vdz1xUCiEt7SQE7fmeoPE7Dz9cttVoO7AJj9RUFtdRBzE
QOzV3xjS7ruxjfrmq+7E9/JLy9QMHGcSdq6IEJk6E2rycGSywTOkeMEyQ/UIFY+E
8KWNIf+paw7uJQgd7wERkZdwhRxLKKMoByWYBQfiEc0t2YmqTkiwUf36Mj2dWA7N
uEMAbAULXwiIK69M4qL7/GYZA1UZ9FSr6rsplPkbq8JQuIefuiWlOienN3uxnqUt
rhDCr8Uiygn8HccKrxgPHz9MAnZQHf94+fRNMIj4ADt3MUrRI8aI5dul3aM2YhJZ
M+njAATfuXTJISCBwMw0IXx/LzvKtpQBHKN1wWG4oXOr+qR80nB+0aH4qmZ6l3PE
py9cX5ydo9N14xa63DaZndyLn59SsTjDWUGiW766NOMiCDEYPb8pTqZSEqX88HoS
XaiVZMFKU6Ewtthx79h1dnAKgWflX33jPYsrmdxlP68l6l7XgZIXuw+d/vTIlOB1
3AVATLM+842LfTVqLCjb7Y5QMtsVlcNsb34cvTTt53aVu3J8GpUI1E0ucuromKk0
KqUHsYDGK13/m9VcuRIGxJW/ZEq/Z/CuhizbBBBAgumEIjOBPkVMtspFOqWvgLbv
W4vB9QbI1JqtNXNN4T/1Kc07ntfX1vexW59lLW1I2KLFClauvZpGv79f48UXYnrI
LhXgPF/pIxQlHySzeCa/o+tyGAgG2UWo0DFFX9utiiDNKg6zZDpGkqzLdP/c02Ef
u/MhApI9rIN3AwIBlB/Y84c8NlUTGQy2DQqUOdCuuPWBeIjDgOY69Ib+2Gz2Ez99
YACqLHnnRsYd0QXA2q4mzwFFUy179dQ3ht3BntONZuhLEgAdz3wl1Ffg05ZKS0Ii
Th1YdpxBfaOZPlit8Z3Jcdvm8F+hivcTRId4iUiVfx7oV1Hqh68xm5nYebVz8fPG
ED3ym1jPIOpWIKrJ6DahfO2Jb+bukGXSGN9DM2nMMTdS19kJTxBsw/Ym+b06BVMe
QknJiN7nuWf2FDk8rL8j/QZBmvJeMr1U37PDIZKUBWuPFdFd7Cad3ZYSrMhTNthE
Sr1mYLuBRrphvs4QL49dbKiR1oXWoAX7jyPSq79075UNlEqQOCz/DgOS7tCvoHYn
ZfalmZcryZUG/kx8RNphb3ctFtntDx0J0jd0/6taony4QV7WNVcep8+QfjltDAQt
QnAuI+8XW4gEe0pQLjE7TWxggzx+sXjR5oX4I02OxqcXhdOjw2erEIikA+3gOPkj
2myZguW25TL3fgx+m7aFsHK+Qg4qoD7+tM4jo2mXqxV4MIjH3TXESNirSykmBfFh
XbMb9UWRhj7HkwyePRR6YAHZ4rct9Si+3EUX9BFtJAN7e70eAc0jxImCdmDzHMAy
w4R/BKGUeM9TpPn5rVxnDY5b5AZJfcWiFWC10+4uSgjXx2IoSz0zQEq0VjWIlSb1
RsIDAweIk6vq64skhxzqaW+tbZrINOdcFo9Og76h2pbF6rXpsFJ+1EWZJMor1I20
wyDel9QSp+QvbZXAwxAtB3QNihWqMqpc0EaqZGA0Hxm2DsZf7g0b7s1nI9jMIFnQ
iLcHeV7uylajvownBlKhI9z8MeQr77d4E/BoJcKCudkxKMF+GTGGn6WOaRkxLhrH
Pz3YS6bsHFXZvgE+ROFS2F9nc8+EZ/Ee8PBvn/Czwrog//WHZCQG7Z2nOhQAljjl
1j0xia/8OvVBQgOnaVnS2coG6BNlWz+rbKTJJpRHrAkw+BC7qboz6nBaLH9/+feL
lxleHfT9lb9B75Dc6DlN/9ZPq+tRCKToeFsGiPg0Oh+d2TeelR4X0zuePZEdOHzM
rnulHYLHwPGIL01v15MwPLSfmRzN37yQmhWns/1zpP259gW5/4vo2Sn5Sf8j6ORl
Fos4FWSX+2zRYXF6q1HwpV4S8M+IKICw3KhX2WQ4OIisBDB6UZn620wookDtrD+J
lYQQCEqGi978SZD5DmCGMtMQWBaKF4zVFHFCNsJ5IwoHSGLu2M4CYuYI3CYJyK3M
rTZn+jWnytZleGZoVVVBcmAmf1zv0KrvrLklybGIaSXM5cCeIM+EBUP2xrocTQzn
zt4ERACc0r1p8hkfbKkirCrqDeTNhalui4oqhKdL7OdhLy89T4xZSR0iLklGqkNF
xJnl9Rk8MOMSMKxioZtFauFvCmqYH07kbIdVg82SaqsvF6VosGFtViLRjS5wuAMF
muakJxrPo6qtftxrTttYtpH2If4oYmclVtUaMSARz4m7ahj8E5YAGCc84gcHhBiJ
B0mqrQllR5SZa45wiu6+HHxKsfMzOgzrdNSYZ1d8S+Wj9CBsfnCZ/VeWjXBXS3pM
omNHNm+Ok1l4CJev9bvKQfXHFLq3EOwZUBGXL8EAp9CtR+xKHYvNCa4H4xO8m071
NtfhpAo7ZQRnI8emp+CIchx/6oqRI/RrfSrG09gPaMqmUuePz4YQPTwFebK4saJ7
J8KPVCTkCJOA3yDn0XswHUAwJPaT3AO+1hxunha0oBp/MRLoPyWaZJR9+k7pwRdR
0uwBK+Fh2q+iNdJ9YRJbmUINh9F+5+NYZolETw5se7rvJ90f79PlbmjaiUbHHJD5
AmNdV585Iw3SU+RcC0iHgCCuXH47r53d3bA9d0qxZtnvLh2Hn3DjjIxui4ESZhfn
ejR5XWMtLF9tRFmS6b6SAph0zW/K2EKgtHEg5bKeQBCX8oYSyQTJEa5V7PBLCQdO
KWHQjEKhV4alpubE9j0h9fO5zveARjxcFimyyi/ab0cv72qDvEJuUoW0yM/Me3rf
ni9SZhsWY8LC6EMAl55m5PSY3xelTPs71dJx+0Q+hrepzsUVTtk7YduZgEny6rN8
QGyOZvtxA40nqV0PN9v//YzplTmcDQ1O/xiZB17/fCb4Tn0J6QjDxq057sMl3QDO
lDFxbRUWWcqpSDghGmCn1FrDFrHrbTka3ApDqshNYil/sggUx5ibWnlOZGv/uw9e
8B6BODHtBxS4nR7ux9aAW06sVE6pfyGGE9PUUkvqrnbQ7wInN1yRGORLPA4DmHPP
EazH0a4OPpHlJrNoZqHlBgl+U/gMq/PlupV7elH0dB/4uYcXmqBGDyjFT5vFmCvO
utLeeThGiG7ibaixbvYmx/10fSqoX44fbnv66us1ndT5o3DNVQF26LOBPWI0fP35
udFKn3oSjZ3O+wJjf7Dod0Bn3EGR9DMKjUxFxppoqNwTIvcOopc/DcHLILPfHmug
ZrW3scaFMHZNEiIEa+KaW9Iz20tLuolzGzDjKx7LaVwaoUuSIx3F/kD/gQHLo0Sq
yySAeUsBFQiT8D9HVOXXjq5ZRXBu3NyyIfhU2tc9kjKY23BIi/5U3R9qprhv6p6A
uNlzdgtOiWThAJSj+NBrX++XKbJO8J6iiwhMKeBtn9Cf0nMM9+QbcplkYDj1CmQX
uonBRX+umDz6VYi3zHPcniuJT05FdfmLVySSwSaEwVWbC42j2F83D+LCsgYPZk4x
f7Vnh4r3Xvvbvz8XxnV33P2NNC/wxdE0a4S6j+hQuqlA+YyNh8SRC9UvsM4k8kzg
lVmbqt08P+N8JlsKaJyiLjrWjmQJrKqkUpw9dyk4gokorGFm26PjfVV7o4rDR9At
8yyk/uRnMkM6mfeX0s+bxkhSdoPiuqWPkpfHtMbfHbQ5bDlDGxLGFir2V1CjDVVA
wD1Mhis1SpLag1rlP1i9bBBqfqNMtj/ZeqrGUtGIxWqh/hCPdCpmuH/ahkdZgYud
4fyGyQ4Tu2k2ZjQMMNjKu1JeJpePDaPo7IPdl3p2GmKezPB3AEcjrwtfKxz8apy3
7um6l149BN9+HP44uFAP6FWDUR++ELj61VdgXBuwA8I6tWu9EHmOkcFDabtN5mwO
k5qO8jA9vf9FHXNdr/BepKro67u3hma5NPgerYkiJxf1WAtEbRcPF4E6kLSmnLbe
ClQiWd1khbxmvRlsxASPMXJFnqIGWcLTc2bN7r/VZH65FpiGas9lokYlqb4fe8aQ
3XCU/549A1Yvbl8I+1/lzaOk+4abDYeoHth8xiP/ehf+VDDBzf630qBqCw+lMDyk
d9UXTNqm3BNmSlstTC55pxytwK8h7He2ZAU3lcP9nrasA313+isL31qTBVZq8qLx
dq8calEL1nPzs2273zkOCg3sZOnJp2kNYwDvuR8HNXH7RUFW5VufNcSWAQnProQR
TtVEw7FJH8GGunfkNlxOzVda9f3oSW+CToACAcp75K0nKbG1w1fc6VBgdhffHQrM
LPSYRP7+gZkZry+SkqJLmf0ltTK7fqb4LbehqhKDlDshgTBazmLvoT6lfKIY5NmE
DPHkSIl5VfbYtquaRQUW18h41q3lg3F4xk+FT+9cwyR1pa97WhMBPRxh+iaiGj7G
EYSiJtyIN4zuV4v8eDUYK3qmeLkHBVc8kZ9/Iktz2TNyiBg/Npz+1vMN9y3x8E+J
gnO83ojzS23dnMzqCXT+sZ9r1C/vqmjBBZpX0uhKGAoItSCUPdi5uzsGNOqhCiHa
TR8bZKCrKLEzmXdnwh8kfXvGDeN0FhIxrd/u+JWcDNNoaKBsDSBJj+GpLaf6zMeG
kWKWEpX+Fe9Dgk5xHPzAKk5Hsic1frFokuuqUvjgBjbCuy0LjP5sPs6i5AQL4Gm/
OQVeyrxZJMfPIkXDYBlgcl+SYVF9nbr6e/E+UNgLyn3E6gFFIw4Z8+145qOWRhFX
H5VURmbmRlsZ9Zp4EkgzJ6gzq6JV/qk/b0tDKlA4IMpS/XcB31nhm6u3YAg5Bs/C
H39m2mgj9RVvi/wMvmcHyj24CIWVoruZcjxUibNRN0Q2+QwuLoNiH/UbxkufBwO0
X0PG5H7qC+3kJa1aU+Y99vcXnb/0WXLka2F6HuEcJQWa5qsofzo2983y3dv/b5JO
EuMZTFnOY3CixC4puANLQNQkF4HtFNPF7ZAUKpliboFwXukTR13sDSx2+2eAl1TQ
MIcbBXHaoGMHjefB9unVCdPWWqgsat/R50lUi6LitvRkvsl4Sd1zQLPrKxtf4WtZ
F18FGZseOYSVyY0IUDCV7j/eV94+dIA2SegpbE79t6zcnuiOoFhHo2OowSYQGJhb
RSrSF9X5i0HiqR0JEcPt7zugKHNDgJdddgTZIAGX9lrTucWOwdsk0NcIcdk9xq43
E+A8Hx38futvKS8hrwD3cdTudy7fk09rOwpcdJ6y5QlVYRhe0xCBrw2qPNGajgC2
bzN52ilaGWUjBbuM3vUStmhwmwVSZuwqWGzMwZnto4Qqlxe7wLf8CE0DfIG/mlZc
wXtNyuKmthdH18WGtwULTAyrqzIEEjmF6MN1N6V1yUWnj5d7wOjci6Jsnkcd51nu
DOqBvfpxW5dI4DilMpZLgf7TlpUoaXKKAlwOrAn4W39NazzXJWTch2nSsKUmlVTK
dmiFrBdtlxyh/HoITYyFOYoyFZcj3t/wOET2cVhdccHEge83Mn3g8OVVbZ0k7O1g
nWvpa8Ukoton8fB35ZVOSKbiAqq0kgk0PVtrPujb0+VlQTiJr9QBEfwlrDU8JkuF
9nwTSIf6wGRF0Og7KoaYXu7oybl7v8UAqjXhAte0GJBa1nn4Pdsy3aneWrndfghV
NHrfdVIdXpcsgF7+zBsJ9nkHFYxdRcfgTvlnQEbf3Kb1uKffh77UayYVhYqYv1C6
rsFFmny+c4sZ6F8KIj0NsgvzPjXa4AaIkxJIJhD/b5O+FKBpMZWRWZm6GOr7zITo
bINDJQAKDs4GDPWqO6RswHF3JeUEOPficS7JIljNRuesN9UvF8fnBAF3v00wS/2K
ZzZu86Puy7ADIE6LVb+GhcD30qKO7xA6HtvjEeXDhOQ6+a8DFC8/x3RaUuYIlW9z
rgtzyrZRQdDxZQD20BVrl7jsHsy2P+RghaVUZ/vDhZx/iNs+sZAoqqqxJNjcD5rc
N6pNh3AV1dwVYtN2R45hSadAjOmtsPLsCGqXzJzxuAsSLW9mb44nhxfH3FJlnGpU
PdcOAXA89PxN6Bk+NlZr5Gz4PkNRqzZcjxhx9oOnvQ6d1r+q1C+O5oX8XcPgJxjR
74mLXKTotxMbSpfgyaztEeb7ZanWg6q4MKW1frlNBslxtXhff0THJU8htCyiVTPk
du9/fQlQLInQZbVQh8DH4c1JHPx4DqTs5sLckACB194gy49BQddFQfvzl4wnljuz
wAijjSVz5AycAgOJA4y7RwMNiyLp3BbtA4w85QaXHiqvJE1BwLjZLQAUiiMifWaI
D4W0YZ0uC0nFicjE0xxIr7yzXo+q7Z6wELkgABwFF6F30dqVUf+79Fo28xDFIpUG
iqsGWyFAFznWrvDys9usYAOhurMW+QFYxIeZIuNpJ80VnI4HxnuVbfptHZl6WvUg
sJraFAw/DnCA3c075G5nNYa4zqck03V8MdfMRG1ZNlooBd+1YZL3lWE70L09Niuy
gXQZGEfw/6xd3fw5F2gxxQPQbM3L/bibK+5o+Vt8+pu8NPO0WlhedTcsHgfpP4Rd
+B/9ET/a3j1LQQOCKAh2CldXSpL4k0JOmwI9e3LeP+5ufEvhHYPD2WRgA5ffHuzU
+52nSybfS+p2G1Z8xQQRzNwrIAcSNN0EGIQi8dc0VUISIsRHxUEAHGC2m0oabZu+
2fIKEnvqCRr19y463L9keLjlccyEAoj6mfxHEuKQO9vCSDdIv/DXbdR/z5s4mrb2
TfmbS3DNdklMRVSkww0C8qKNi8YADr0ogdeRoSeFqYxb1AG13Thoi8qgyP+T+Tsr
2JdcV14kSodTJTJckKxz1ozpdnd0vhKRnqIIAfCgvoTSYQLmuaxXg8Ni8oY2g0o4
gkg+WD5oa4JDrggFthryJr/UwvGt41Cf7bHo1UWWcE5Ut7Jdr6ldwi/LMPd0zC0V
C15Qp9smxqCnMohY/v6ZruZ3H9v7UU9Lw5T49VYPfkUPk4pN0kMF8Hc81zoehAyY
P/8pmhDeGxwLFj4TM7zxNc6MnYzEdgHZy47obqocAnyOet/klqmmhAtOElPnRPbs
Fl/v0p78prtn9lyxN9wgLe51aZdoQUWtVSAZxu/ioT7S4S/4Z572BmdlBh8MRXQ7
4Hng0hXdKBH05MsuIAWpv8lkU/9/XgfFcgBBjHgaD75VJzdQvjkIMecZK1pi4Tg4
wzdFn0c2c4ScU4D0HsZbkgDl/eCSF5+RoVpgjns/951MVjZctsFpgKTLGpbo6Gaq
a6MDyfJvafq6mP87Vr87u8/nVVZ0F/ekdAJLn6Iy+vpOVQDvCaicbQ7Io27d+FYY
Yebnqy7i1ZUhSXi8BQnes0gVIHn9SMnJG4tLItRIQv1ina8DLby4Ohudg9AamS58
u1kI/UPuU2e0g0EvSdXVKo1+efBsqtbdpeQFBGdIz+VxN1L2ohHeiHR1Q3+NMCeC
Xq8LApcE/ZQUB4RjyxvGArLiL6vtXMpopx2mvLOAds0ytpGllTYvSm7DE0GDI2gW
+ljPabK8RGi01JbqeuYViFeLG+LEBKk9jf2HMrxKWWO2Q7mmbkOe51kQzjNnoPoY
i7o7sm5NHP+NYcUieJKY87EdKsbjO51km9lunQ3zdSyq4Zz0F7onnsm9L7Tau8nO
NT1qBlsZQsSTQrZQTxVpF+ulyTME8eh1qI9h+cs8ivH2Q+B7o9PNMCY95cW4XMi/
YSTgT4+w1dtdo6cQ6EAqs/eiREMAAdfG/wb05XbglBfpbxmBEZatqqQ/ggwvFbgM
QDqbOBnIhacFyLccTCtLmadqpcuMwpcmKhb6WRDouZgn9fXLIL66s2naYGCuDMiG
HfIb/62bhtawijXct+8HvORXqCBTBIRx2vgR/eZfsY+KSra5UOdyogPBGdEqhnPb
dT8dzkymGUZIa+XdHFw+IS06MC7KaRAft1LLgexvqJH3rBdgYpOpv+bYgKG/EWpT
oKiXWhtPMIkmBOpQCPWUnujSxnyCFQdryBImKZRnd0UY+Fil7xFKKLHCnsc71CWR
4K/qofe62c4WUi5GMfNsYS03ovpXKtVhZvWHXXmIYeG22Lhqe64wAMPrJtpND56j
1MIymxFX5tL7E/gLYOnewQ6tU7Xj/ZBttQbnOzpLUPXceQAEXIxWJN+fLwOgZlt3
DmtlAHXntnmUe5nEzp7Aae3Qc4JEu6crrwNbd5otraTCc4qOuSgLgL+YBbgtxEQS
VNhPXR/x/hZNNwLV/t2xFvYkVuila7Fo+EC9fnzCuiSd7NuA/tTCddSYRLvS+9iC
i8TaiPCyeue5zD1bo0CPptP0D9JkAp2VogHPwJC68AirE2yO0nTxiDrCVPHW7Syr
E+aCgLqxAm8GUkPK5vzcMPiLJXb56viyaDRUTB046zjQaFKcg3WtviFemV719s8H
edp5l7gDyfHOD3VYZ75jr/xcLT0/DkCv5aHvxYkF9nFRGLPSk62wD6xTPRXVwEUF
uazpmYp4YihnERJNwCW+4XCh3V5OIstBcpG1TI3kEYTQ2cOdDNS8DAY7i41dduFH
tRtvQGzMHWOQ5JEfuq5Id59PMwmp3pQx8aGHa8VPp9xrvq7OL7RoRXREHuYSs2LB
7WIj4Omj0Es79J/qGCsXL8ub0TdZMfZEBtOk1T129RQ4jnU0U52kpcQ27T0yK7ff
BQ7cv/C2K68K2TtNGVxFMvqPkCSPzxRQhFcwuWhbLgDDGww2R5VTd3liiFnjFXQq
S4irm+YoR9j3tHEr7z+6RvQ9YIUF9psXvcAkW7HUbVqoJtHBtRxqMpQjuosbkclw
tt2y9D4U9wZbuxrfPvhqpXxX6m7CDk9XSQMAjXMgNWzIbkaPCJ/Io/ZYWowvdU6x
t1+kqBVeMidq4j28eeCFBXZpJYmUZVtDMBpSpY/b5RBh5adV9fdz/t+nMdEY7sW1
R8un8tRP3dDH6irA8z9MjySoA5KZrPMJkGDrLPqxCOyn6ybx0H4Y/HvLKX0po+b+
HBSwzfWJ6FoIjPa21TJLeLKoy50i8NVVQzA9EaHwYiiBxh44wFbV0h73XeQRxx55
S69PzDLacGEQFB3dteaZdXhD3JWgZL1j7SzveNBLpzc140zBu0iN/wACKSsc+uEy
S3eWp++7a15R8rFYN5v+X/ujgqHMg2aT0YKuZgEGUrNliJpg+rmlcJ0J7WzFsYBB
cPW8WXfHNnH5BWXuXwCty4zPU81nqOnJ1/CC15OKHPmU1m0VAjlqPj86W3MPF14B
RPg09eoWYc/8u4fsXqJcAgwaXx/8UA4GOQoIHPlsEtrRH6ktOkUSVZwzbqtp/hOw
22q0QaZ9i9Bqfk4jwxmC/H+0Qp4pgawXf3z7LPIppqBy4BxzKkQqE0bfvsJEPPEs
e2S+b1Iaouj1rQEKYrDzQDzWjyj1a5KaYZS34gsqRWTZDgXc8ESWmYRd0+QQamuq
Rex5m9/8KlrBtaC4rYmlczdzVrk32qdFWvMhLxYAqalvLRnRq4P3RIueBmXXZjLM
TClAP+w8ZHbhtfYUi6hEWF08+Aue7ZDAT8bwVx1ieV/j57aHhl49n9Ku+H+Nd6g0
FzzIHxd94kpb4RrZkqzZcpXVOQRxisGLUSCMM8FRVZJgHSNSM3tcDriUoAoyWwyN
30WVgeOr5s+dpB32D3IW1yyatK5i5AlIENFj6heePRnk/ZQ6NkoTWsiLnAzZv0AK
FyfGKwQDDd2OIQhSfKUKhB4suwa6/9lAdKtf542W6KiXfbvATf5dAVwBlVfZUQFl
lOac/PgJaZB2CrvhfpW8gaHm59QXo1EsTEzgTXfk4XAZUjAeu5LRiSL94XchQlel
3I+MBLsdJR6ChC2XJ1y80yXk5I3wd4BO/PletGWKUQnf28qm84It0o7HhIzVw7Gl
moO7dowvKG6Ahq/tEqwq66bS9r8SbRjU69L348jsduJmBAWRXqQjEwDNI/F36aeL
fDSsaxZvsWisT2F0NZqNWz//6V1AmAFtuh8JrjB9R1Vax6L7qc4gLK02oQavA32M
cJUZgoOP59dY3jyH3KXz0on1kjTF00DGkcLbqo3qqSn1Lt24NooYLd+2PRmFQZGU
VAHFYo/wxF2Ly71uRB16/prDvzOiMF1TZ9NcLs0g4hrtsm9A6hsp0Bj63Aj694e/
ZKfZwFt4Mt3rFHqQgzxRvxFTBNS+atW4Zqs71ZNkx6zolVma/zQYvxtGF8yW7pek
L3D37YQrTPFdXjz5bVkiowgXjYJyDhahWML8jDSPRUq16bFg5IlrbCIKuTk1reCb
dSohwM7ZcCdD/HvMfCjEhuCJzvJxqxXpz98z2ntNK49xcT+KuakWTTgEfsp2QLvl
l6uAgM4o4m/BjE9JsOqyKj4V/gBSHePRG22Ng8jfHiUf28TCsbPJbXJ0TKXVlS/S
BY7f4MPGibHiYGN17V7ovTYubNtj/Sz+o26BUmOSvpaKr/cPoYmKbLfnPJU0iKrR
8k6WhHtSjKUoS0Xg662Ni7yHtfKZMC5E/g8b2gfY7/e9NWRBVHoYoXL8QCeyFnMe
j7CCm+Dwz3PhAnk7UHOSFe3gTzdPppnB+WiNEedTfJzXG6/+A4Lp3PQoBVKER6+b
YHa1+ohAV2vs1MdCECUjZzg3jBQw/D88/wZUMsyzR6Pa3x9E1w8PkH2bcE5Ngqb2
h3zp1aDp3SPUuYWBSQOlRHehWvXVjbCvosPjEwS1onNC8MJbYnDlOV6b0s1kOogp
x4xn2X6p2vImnojn8NWY+qDiuw1eDKpPQbk2ag0A6gXP7DcNy/Uu1KzDwIvsZYZp
8X3KlwLzj2KAYgNd4KtLL+nIBBMIvI1MzjFfez+7GbAGXwTjqIhTxDKg7DKOIjkr
LIGCSWe4Kt5ocC0eoIiGrXECsIm05ddZSUSBD3J5PwASXPaI7hH68Rv1XpM3K63S
TRHQ1fmBV8y4pJquBYJDmLBCEkf04UzR8ULefB2Jo2k9QQXUCagOHLOT+ZdJSWNw
brLIYbzojgrZlQc8kbq7uY8nWlz1WTBUWD9JZPBUfoj4DOMsRlzJZDGvAG5xiz0L
mcAXdLznmtBHlG0YdxBcqwmWNam0huDbMRjwpzYsY2heBTpyKosZ6bFE9PDCbfnR
Vyhacx8e6eRiDX6mqNYnomJ7WUCuUyL1whLcOcZOPU/WwWX+8n48brNBomsfTPm8
djfb7Sg7B0JFGZTAltV+r/GlWlV30UIVdpnKClhOulknikmHVUmXuTxaBtBfQpAw
O8F7Y3LbS13RD9SCuE/qidFcYjTz6SDPfEuZK+5BREkARS/6pjOtdqUR+mUSyhtU
qLsdo4b3MDXd85YCZLWT1Nma/mDOD4s6omf0flj6+j6XErNYuUnSAdqUQRCoJlrf
91ZsjLx6w3C5dCaRwn5RhalN48+DIx7tMf63koJdSjkkLIa/FAaoi1GFAhlrxpNK
2MOGGccfRZMtgsthBlzHTc3Lu9sjLkxHxCv+SNvTt0/xC7zKJVsNRv+tnv2VOsXY
hFV5735x386W7Fy9tvDhyRvpw3b2CgF+0KOkw1CXJpv3oNhFr6oSo5UVlfFHMfKN
duhPOcg0CsBn44pY7Rci7Q3JfvuEdb7N9nJjMME7oN/S8s9VTStEhuB7VH4RLXVG
VmO0xjTQbhcG1pTL++6H5yG96KF/kWnMs5VSgFmEm6LX5scfAUT2SscN0sTW8jWo
LExqiRyFrVivh6SBkxRTtsLQ7UpQVrS4m6E5xFpbF9p3Gd1Zdl0z4OzHfSNNIU3r
LugUHZtStAKDlowTljgEsWFm/+nSoIjA978TOXSpzAK6Xgvawj2TJHXxU1XrLqER
l3QkV3t2yDxmTVSmaZMYoDdR0I0UX1IpgQrLmgqKwFeoYddRwdxJ5NReOI9WhSKe
bgZs2wiRoatBcHCyuxXoimzQ5WccsK9lv4aIQIMZ10IW+URQ1XJdj5H+1EVU4120
da+RyMnD1SFYNuiaDAn/nwsvZMAlGi7tjWIj7IBILchoEm1SRj6ZhkP37Dhzkg+g
35jc9X0gJrUBlqUPN3ov+62PJ2xeBZvEBZDJXY26jDPXLSKwgeQxkLEN/Orio55v
jZKTzowOhN0WLgsl3u6idIovH1TE6ThZpx4XF4EIuo2Ms87aUU/Vg59xL5AiDmsL
k/+lbZyJs0khkdW8bjR3kTKU6cwF+TZNDZE15I6p21R2V9paiH5Fl05mmW25IEo4
wCAnfBkDFa89GL2CBqM2Zj+tcFE47EcwRM1FOQYSDgodS8XNDzW6TNIbMtYkpoW2
pJTUnoq5CYZF7FJuuBKeaZeh2pgqnDkrPh5WSVqqABDjFA/8m5FT4wC1vh2xrRzi
gnhhY/Mm3QURpI+kxnC+FVH1P0AQQvjFtaPZ9vN1YGfdwhwCKJOCsHyjQ9y+/AyM
VaxIqqH9CuWdxigx7w8azpbySfNL+W+tkjW2uaMSCnfDtowbO+eh5vYQWZMGgrfR
R3RjIhQYZK7pxQbVSWe43zKQyhLFgoE+mmwnj/gJeZ4/hFpNkJ6XF9mFnk6uiRwo
CBtD947hUqPumYX/lQpcMzb48GOtL41Fw3oBTKJpMvgbUvgZh1bcFPIytU7Y+lQS
lJ0uvv294FG0FnzE59GzFweLuJUBB4MfrBrhElzCDvb0g2UU54xfiZb7qRinDCuj
Btq/uD4yacaMidGcpCE/l/WyB4YOZcCsOtrfI/JMvIgeEBn7XnKBiZ+gTwA8lAxC
KqnsqYmSaCxoCIrrddfljYFB8HCYjHNTFGU2o0BB+UL8GZL1jqAc2K4TZZUSUzBW
7m3ZrrSk+m0voN6uEl4WMNNh+7GLPkL40RhxfCkIsAyDZ92cCWMEhsrca1etMbAu
ZSuBKhh4O59Zu1aCnfwowZrofnYbKejRPJ7Ad/c0PZuBxORUROjGWkEK3IpIbCnl
joGEtfDwpluJn3Q2UaBwA3Ai/yLwTbcgcdzINDSsDrwPBObfXriOfrPWwQ9ChfwL
I5plT75/Yig0sKJksyvHfm+MGkDzvmMK/PO4LSS8sMZo9Gm1qZ8yBhwWHMpuyHF1
3tjWiTmWV/BHviBlquBz90878O7zVGYxV6+PwIgbw+JLs1Rdk2VR/FAFaQgOUNTB
QuAEJ0OlreTF0e37kxDPny7VKLDDVyP3ZpSVMUBIAbdDobj6iG9LfiOpMhc+22i+
vLa7tcZdOp5rQ34X0WiJrwxTiQp8haizG62C+FbXSaoJ3lEt9/ApbY4TU5FUSIZX
COBnFOpCvgfPETu6OBOIuSTKXy7bM8PztO6atfon1uuvWy6SBH0/TrDcsMZ24eNt
OkDeJADPdXm2acgqZwR7BWnQoioI1TJyAb3anziC3IZkac4rF5I/4xbWccPv8ZrZ
P8vy6o6XE+Y6OQX6XcXH1dVcuhw0fZCd/lGrJXW1oiTm9Wc2I85Lkb7xK/RPvr7s
7yDwzR387F1l7nNcwk60rbz8avf2JCwn+TEpj1Ve9UMwCI/Y+UXRVz2gYMRt6iRM
7yxKDNFpOQ1lJsurT9KP8vR4Vp0t84fsE53lUtLkHRi+G2zTtMcEHWCxoNtkZD09
URmCGsbvCnwzhNn12ZWMtE0Hct+z+Uq0ImfoDQykFcnyq41XJgZ6o1dBF6U5/6dk
zg3maX+5/yLcdfTCfUDs4b/R4QxIK4d7IEJ6BrY1x2/RjYsQ3LTgfcJkdyBwEQwt
wkAvwDuV+LQNbPbcNQjgaVM/k+m882iXZGzyu/mAchtuJHjiX2GFxx2IYiw9UdPi
tOXw1rB4lBGJy26tbSz3pJ3AJ2qWk99MMUnuNbCXrgONBE+vB4OBa+7l9UEyFIjX
52vvpgGRasCXJSG5H7JQfGcbnOEqr+fr2OH+5vjGJ0CBy5sQGbhCqdDmTIcO5Qui
7+oCGO9hnL6i2yR0RMRo60uNrEsEe4EjNEuqDhlb9a6W3z/dvXrQUPsP0PHwhYzf
9kkHTY3GqgvuI+qSXTNyVAd102SNAIex3pv1T91yMxoWn0VHi/SvXKuE3FxlxggN
T4C3EKoo79P+vluqO/gylunC3jqjaC7VpWUjue1bgA2k/IsabVPAUv5bsmFwsgye
PGEZ8We82fnoA7IXAMPrZd2HrWWUlidjKDP29RJvrO9DxA5M15MRe0GTcd1FJHNy
auwcirYLafXT+xhk3Jql0gQuLQppt3cCwzQ3GAfHPVk9PdA5CynynDltnLHeghCh
V03rJbVTCaIXqSyf3r6exUKjkmXoMiXm731PFhrZASbW3svn9/2tQrycPvBxBy8S
GepiTq6pLOGWNP8kI7zBtJTzHc5KINfiqDW6cbEB8sTEHG99nHJ2QqcenEaSHMXb
2NVep6e3ipMQayNrZ0AcWBKXryFq9xUpgg6Bxuo69Mfl5ie/xxvTYYn6v+8rAF8b
wbRW3YKkWz3qGipOTpU5YwaPgA8O7AER+OJhUJDy6Vda3cVnSLYw2qT/u5o+8fp2
VxHxHpL3Vkx8TAR5/RYjj3KXO/957/CfEGkxbcF/o6xUZC+AArqdTijQYrwgxf8x
5jed+TBijN5GkHSp7NYdU6L9/l91NGXNeDdzU01VamWksiKhgs/mDDQq2Zul/i+h
XQt/Z8X2kl1rvOibYKqd0iHTt4Unp+v2aH1gFJljxRheY3N3ifHZ9+1fK3lfES3T
6pSef84bsb4f/2laLlaofPM46KaHoTJ0c/VJiwLZ0+gS4cKxJmkhMznuzRgcrI0c
wA/ta9VnEU+9QnC3d1/RZWqARCemD7vBsfFdsMyaTZ3ePyDXmfQ9C/yR4oz8AZh3
x8qXswSxuHafOl/irUc8Y6tO0mtBERTzvUuCGHnamsOMnDnq0LiLYQgNBaxrO+Ll
4Sxa28jXP7UXh1jLoyYI9uoTsd+Q29O8c8hXFBP/4sRR2Ugx8Zi3CHwMTqCn46Vr
1ULzC38S9ji1yppywanzGYBuLQ2zChdqWKbshkJBQP3Quai+CA6vX5ccqH48YIsx
ORgmtVZpfQMsclgfp3iSpV7K/TpTg951i8qUGvzifMFiMCszyMnjEob93MFPPVdv
yr8Kw2CDiIEeVA9cCb284Wow2iLuCDk988Aw4ha6kRHkwt9Oz5Y7CF//xGQMoaP0
ZBeoGzFVj2p+V3AGJbA+8zSCKKaGLeNVp+iZ5PAaHVpE4CMbUir0GFvYuLZg4xls
lgXdIvV+ylML2AYu2HoxWaVseNJvbNLyOm88vGgKrsFrMI1EPi/TxRvKYBfBkDS8
OxVYRpcBHyONqM7SlF2o72lw7VPnseDeyDIwZ/DSjlomGgIPLnml+0U8J3bRdW49
C6XNmgOUWcrGk2z3atyIOAV52CaPrPuwQildNMAq0ZP8+OrylzEdbGViEXszmMPj
Ra9zfqEGdjPUoxBbr4GGXPnj9T+iELnts2Yi8FIsuNHF4/cALmrtvitQAqP/Wf8r
3TcJDz7DzO1IoI51NQF5x5cY1KDwgEjQbPKlmvpqRyRwtjS9bJRw1Hybf5YeseFd
ZH4MLyGQt3HoK1FiFMgeH9H4VBpLY5HZpV/WO9HS33UenZKs5WfDQ15iBKzs1YGp
kskX2YMIJNUgEKZEWiaolh8gQ2LFT6eDnSrCBBLQ2QVE3eY9kX+4NonH5epfYVPU
E81VG8AGZkhEFSQCSovehsiFj002X1DFJllrQkWztnp4eD+l8vHuDZQ8eV6s0iVR
0zQR6vmbD/f23q4A7FPHlFhv8Z08FNjd/k5PWYlG2Dslzv5zGcwmt9Dgpdwv+RU4
h6nuYWCQoznL9s3Rjn8DVXm2N/0mnVKdFAE+D1LMoLFsWai1zqBakwwfCRc3VwP5
LeIKd1j5zQiAwveWV/jAgYKaBELVzx9zDNzGtPm7Lag4Gzq9RWlGz0otoUHsEGbU
wKYTM4/DgOAUnHBAx7/gDUFI9quSnD0fNMAyUUI67wTljFNTHjJ6C3E5e5nPwjHk
gmipJs9CczUHEXgp0K9qofKB+N9xLDjXywNIS0ztBmQtORBW8it7PuertFPM3ntg
UtrKFGE8kM8XLgZsKGdZAzAMMdICoEze7sMWcPVepNYGSSQYfjCvVU64xCZ4tBgG
i7f3q0zR+CM+5VO5yok47EygmMvZiJqBhq26HkzA5DW7zF3mgb2DMxv66SOSX+BX
YTFjBzOKZlkw35K/QFLtrlkP++HywPnijAC4jbydq/DbtpTu1sU7KT5OXDvqbn0W
S5AfsQSgenxIbyWubsmZ9Pb1hxj8NBvnFwU/2iw+FtmapNV2JbilCQb05sF/ovU5
C7RIAFcKnuSMI38W8UYYkAF3YP7wKI7ovc3Je78JyYYTEj9KZ+W/NKjCiFmy31Lx
3KWi7IRkcZLqA14F0192kJPy8qE5wifYhJ9RI1yEZqnQwYNiNPCf+19yD7samWZq
j7nu/VPypjI4e4Ih7TtaGSWJnzh/KkDCFu2OVzIGc2N/YU6vEdpaoKDS/+hluFuu
bq35yjAICTdPUlcfxMhv961oePimwXYtCTK3kTRec29/wJ/9nqPRpDqg4MoykiHl
Tkmn3d0m90OHp9c9hZ7T6Tpq233LZmE9eA91lWbYF77UcXycUzpw9i/zrVLWnTw+
tqhuKh7NKdkjE8wTgXjvqeKfoYEh9vSN3i9qxU7ARlukygK1FOOrHKL2gxqpnMF9
5BSyPAnvvf2z3fIt7DBY1uUrwV99Ia6ofvW9QmgzQv621YzkZP3XtuETv4wsAsfH
UV3qLK5B08HJZuCtTZLMvrXaojHsb3QQIjWxSjq6WNZM+O5PnpPdpkj10kLz6Pas
HLzzRjzousBhW0uSKXdCLLygyh8jIsbKDeQRs9cwdTnJ5LY3dzszgmxOXg5penVG
AwZDCMB2P+0JYkmaWq28X77EOocyg2VWoRftaJq4VjBxUF7VOXrh19N9r5zFzkMT
abWBd2HfqwWHLR+llZoqoOkwwJAqLp4nNXXiPZDECUAJYrdb2+YjqwG3jHvbhZ8s
y8jO+ViArUjbNOVpmBc/ipYJmo04gl9ucbnSeCbfK1cG/h6sEIz2Zxi9h6RR6WMQ
scSWSXH8eP9FwSR5KhiVgGBr18ZZksOH19T874CeJ3oJ9GZBLqgoU/shIuO+rTNF
93cFkW0RV1RZNxNNcH7ihEDSIt6j/hHTuSJvTbPapaJZvdT0/P6/RZK6hK5+oZg6
GUm9cSnlmHjZ1Nt/fHb+CR+Qqp/rBhygGGe3/2GDoYL2d1q2gO+8l0vGbBw5f8kv
/CzY7i3Kf+ePOhccpg+zW1nCZn8gJpDamPLlI8Tu6YXQv5fosUXTPSmWjouLNeKf
MqRYKFChTjl4rsoDSe9+XUOVkoBtn2Ivc7An9Xmkcs5c/D/lW3FUdKl5qhbKo+ZE
poTSnEklSjtiaAXUD6p91PRqc0+SOvRsbA3hoJXGzixDNsphKwY+QvKLExwb9E6K
H+ZooytlqzC5Kbyz1HOZ/dn4QTN44hjUqnnxfUzan8DCh+Y6hcgJMb/BkpwpfRNc
DfCJyAMki6V4t55rky38FmVFKafQqZ5Wx6kUq0ovxpEvIzqusiQEQXmGWdYZinPE
Ys24LFE6a8mnTsE2hxtIZEI7kcC2LqlHImOMum2WxBZIE+p+0kdNCLSNdPxQFRc+
vHqmt4ZJnVXNv8/hKKXkupw3a7NCdYIJexCMC1+gDxMT2xtNnUfSlgRJaFDBYVKZ
bGbbh+KQ60tB6Rgr5mfDMjgRPpirzfmOQ7ENQEgmmKBfVQuj3p5A8qhLWwZt+h96
vJd32R8moVuIrRRH9q+g1vTKrqQ0a6ZRv7+8JIIznbNRTbz05UyLCsnmQg5OWHDP
L1Sh9vpQjCiL6J9Q/lxxirje9FLS3oIFuIKDlFRKJfBmkVNyjlxHFWdaFsRtJFpD
+v5uiKct3Pv7GJ6gvhJiSr+tpyHdPdjijMEzBPgZlwru4T0goaxd3DW+KBM3Ud+r
jyQs21sWg3R/TkARZU76QSW+1lZhBJ8UgojLxC6rv10=
`pragma protect end_protected
