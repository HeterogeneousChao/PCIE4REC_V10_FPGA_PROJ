// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:15 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h2fqdw4XEcpYiQjrrQf7psME0raTyh/mmCirCUdBD6O4LP7FfICGaXn/AX2TSDh9
eRZLEyp5ALHPdsU3FYBDCo70CHWNNIU3HCKQTV2EP3U5VHRAnvajTtjV+mHpsJu0
C84BaQKagcKeBJkzAN7juXASP1RAIzb4vBbzWPgOFTA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
r77zunKkNv79AM3Jluankgt2zyVKFG330+2PZXGFYC+ukTQGnSmcAXRt96tZw2y+
0RvvJrUxYlfWU4thHmO3Iaa35hK5SSTrUd54UzfKc+GeOQqf04Zuph4q+yEYEcJ7
N5+yqcyBkHFcecWSw7c6x95STdpUCNfTMCSo1iETfnIS7Z9WzYkvd1NDQjrT+6kr
Uszo6fvQSb0EuDSN3/ZIdd+mgCy1ZwtvxAmtT0NZNU9GJWsqEt/aBd+fTiFOb312
C4fLVR/f71flmC/wrO/XkpX7+a+B8mnJ1HnYgdqjJcAZLA+rgAdnaCfiLlS3BCFh
kZa/ixuK3n2IshpHriceDk3plcKeXR5OUS6sjthTpKlw6eavpZBkTAqX3MtXachO
VD+Z2DPmUNoSqt1EIV9q+vi25RkAasPtJqDX+lhpSobflRVEhR/sjJjYDEnlo3p3
Mwh+44dkOdPOVczvaTv6CU7ntANhjBxKIRLs71YThHZS1TlkcqmNvLOkkvkcrzlD
xjvH494Mhg4d+ULnRmP7XhUlJn/peF3wLmZZn94Jh788/bhpBzcM3OdBBI0Hij+V
reoMsOAyrd2/vbB9u9XLOFwaPhwxTE9oGdeFrkzMzgGYwSNesyYoqrZb2sqUtMkI
TcN5+F8aLzWXNK3eiePnvOSgDed53Xoz8WfjCkRxjcScW6UAOUNlYw04DLI1Hqdi
vBc77HwgcCmp5v42tuPIrXFu2JdNZOxpZXXteHDEPYjU3xUsKqi6sEH7/kEsbhir
jm+j4Yr2iD0+T8kMsH2EW0kVKMM01qOmE4f8B/ekqmPwUt7yiQr14Wmc+rTarEcJ
sCFAtevmtpINLlb5wQ0/vFzE8aZZtgKN81Mjwc3eG9b3MMyVB+kbEbXFd6M8PIKl
1ywOMJVvXakavV0cUxNPVPTbpVQBLn89ijEnX/KxDhH0z2PIAKoR+ZJGfsSPzT1y
GtuLe9Mqadold1i1so0A4RO8ff504bqFQR3xF1Ghi9dq4pqKlMHht4WNXb3JQGHW
ZqodOLbW7IvRuXgGujXiFL7wAUVDfVL0YTxMeAbDp9XH15p5YOWuSXPP8dmeydvl
ExgLyrK8f6SLyGYCccHzDheAK0YMSlRk0rwQyyeF26LVs6PLTge3Ht3O3ydtjphQ
XrrJc/KZkMPBIMbmqpnnOgHyh545B3kOqFSEzuikeLYyE5Tx4SCn0GdJ/1ikZvmY
TF+3IYK2+sscdTEtQVVLWpsrmcFFW13xpL6Of/3gTF10MASBRBw6LnvnzOP9tAIU
v5G5hOGnKdAq86MYQ088V1qvpJtPR5O7mr3H8TJ4hFLJ72MfLy04XX82oIRutyEb
/QY7y0RDdMgmTrRU20tuY4QDMBXG7Ir5QtCigXTxfmWAl+oOw0g5E3EA8kyIJagT
ao7YwnAU7es+Bh98P3hUmZw1uwsSlzZWYapoVEBDqV+3n20YrfwHGhug3jpzvXg7
AtansiZKGFUluCTMDfyyfM/aCb8MdJsAgh/cGDJSJOldCl88qF8PCJF+LClJVSPC
a0eH0XPYWYQ3L1302YCNeYKHavRkU4gMPj8rEEfSjVOwLf5UtrQT/4wDljwLY/oF
lGxzKPktz2q0KUIfUvWC28lS5dadniRusHnce4tozYB0787JxT1QEARuCKIcyeEd
t2WcJmGzvFtY2GKH53Cs4smBUrbSpWHXUbdQFJ4dX8sWH/3B6Zy+YoOGX9DSfvYP
MHuWG5d/y/NFV6FGsMe3KmB6/7CMfHOVf7gy2HhdWBg4FRx1TGop4gTXf2O9PVd0
WeRAN0D9jNd5sn8lZNYkXm4KEyk77/MIvTuARU4FIAycaHfpnPhpl4qMUM9V6s4O
yXlcQEjN4sI1pgLOD+I58K6E34ZqOkVRkYN8IsAkJfW/Mjq5zevlmOlWZcxE1P6S
672317FzBOaavvwOp/5WPbd8FWFkcSSa0SK3yWNyN0KE2pppNLB7nq7H6QI/Ataa
TgFFrazRJJHveOeq3m6MaaPtRD8YoC6LPYX1baBl4rHv5FlK+2shtHdqTUJZ9XCm
1pnwEDA3OoZtJCG5Wh5Hzlgz10FiQ9AYrppPp9/ZfGGb1viwDDwH2SW/JLHgi8nP
SAJpG7q7q8lft+lq1i56pQLHcaOkmUtpzDXV9lC8SchIpVWF5vf51Nvp9nOuqAPl
udVRKtpAhX0DnxPGRIztBd5fiU33EFWKOMJyZYfMSahxc2XGOp2IET7Xvjt+AjEb
6inQ9Q4F+cC1Bz0480BXMdATb95eCsZzdgi+HD3UYbE599AaysenqCJy+l3P7hLQ
XZ301L+0q19/1QqKNWGO6blVndWVqXlnONY6CjF0IVrdR4Yi7KvtotYF133+wR55
PnK1ltACOOymNCtwBjaFG3oLiBxXrb9vzTD9qrDFs6wp4RJobay7Jo7CAQLlgWC1
BUKNqZ+e+w++cWN0cKzrWaTHWzBue/AITZzssHkVx1iY+cyFyysWSZMqjNooFfov
sQWQcsTeLfQ6wGxc1rqYnpMmKvACVpKrSgnyOua5JFeRO+cxcR/fPRpfWYfKDO6O
eXhxqkO8CZmZHzsy8EsrddvsevdMwlpSy1wOMBqjfVxi36fzoTVUKRFHveXz+Xa0
o04q8VhyFwgj+Nkbp1s0wpMwiABJb47MbzvH4OsU7A/9z9mQAlRcTZ7M8+j7VJjg
w+rvD/wVP8O1UlDILvnmKQDpOBbSLLQg48XeCjopATxJoYrCEC/GOWWA+jPnjszb
vKQzbIIROwV5zJvApW6QQThqrUsycOpjo0c/FKJhGi5chYgyJbsvpEQGaewFGj9k
qhe13pVa0jwXmNQvl6YZLKcOmYUEqTTad3OqB+x5w2nunahpOgxxBi+qFRI1bnZ7
Uzr0eTF44gbh7PJtTpME/KKTLFMr4MuUCwsdUfQ8UYUt11ae5zslvrlO9wiHrL3i
Jz/WSM9fVnKC+nMqIZQTAywD6ucYeaGvSGYXc45Asjkm7QUdoxmR1wtqWoUs74s4
xWUipnepi9Vaguj1Ut8kBjgATLTTHjlhY1tds25XCEGTuVcDqahpBePbYQf6QyMN
x4kAwSd6S2VhjLI9xe1LEj8VbhHpiI394/n3vSGgO9kCgGCPMerrlZyBqB2IKZ/6
mU/MhOtOXWgUPBWeW+4AQblE5xetjSGy4o1QUnATgrwVv7KU+lUPc9griYWPHHZk
wPkmdVc3Duclg79O251ii2HVl8Zcd26/Wqn4rOgLlYKSZUfXMTOQsYhhz/5Ex3DK
1BLXsI8U0Br53eqxk2k8gZJA8g/9uXjQEPu/9giTKglIxCIoUdAqW8hKGsun8/+o
Dx2k9oZSmh4u7jRsloLPhKKxZNrfmqCKj2TMjqX2jBz1FZI8CBFs94pUrMDt/yfw
mXE8f2/ziF4XJvWjkwZW4F4yhBOX+pUYfP2ZhYLOQPVjo71kfXhOyWnANE8DN8+R
v6JFvijf6kEfCo02FzYvKzUtXowy2+2NDG1NW8C1ympVh+R0DYmDgMc4dOYdQbUx
LufqcLI8vro23XjqFGAGwMZkMQbAPNFcyt0Q4IiAaSIdRF2g2Y4e1tDvFYMjBbNT
H3p6jxlFIKo5MvAhQHfzAb/e5jZh5v8LsXrFvLrN4U4k9J9dv5WEn1hSzpHDeqXa
+1pERXp/7Bi0dJ7a/NzoLm1ot0X94mtE542iv53luixNLSWkoqZSUGzymGQkyM/3
nX3tDTTL083j6slN334fbXz+vfAVqg5gmNbRP+Y4V8bOXeTF8b/59tLFI29QZMdc
/ei2827JwOyLWLmx4AAYdEcpffkFLZ22BA81IgpAXemwsNO3NbeTkCtICTseINHO
ej4Qcfi2EV+X/aw9r36V2DFNbEMDfGVckvnoR2yGYi2lhcTpCOt4EUT5LdoYsrE9
g7lSCuaFKGzGHMV2Bxl9UZUbf82YzxeVffiSz2kT17bCszqn2uPYGrD7EJCtoonW
LvxXgRDsfUftjKPyxwwmRITqMPchU+lZgiIBGYs35FhVpJ4IGnsQtjO5WTzYNHwy
5Z7Ui8Pyis2rsXV8YCdCZ1Zycfp6WqxtJN3eWIYzMTEqhOAZDcksoRV9Un0MInqZ
NhG+HLA4Cd3GZOMhZNgOnusd+DmgsA1wvtTD28E9Qjd6xNv/x8XKmdo8l3g4s5Fe
81WRuwWHIcdJy6ufpaA8iCsdXXj1ifzK46Gvg0KteoIZyX4wRIsAC2DjEP+4O6of
nbLIhK6+kfJH+naaRgoMZ2zfeJf6ZtoIecpPJK9jy4Sd9Xk/8LQVz7gP74Q0XdJs
hXMCsG9CvoXuZDTJD6QZ/I+F1MzmbkHJhdlXBCsJCSxPYReWofkKdLGX7AlnuilE
qW6ZnKy0Bb4eo2JdDadIkTo7/IwAX2Nll2Mw5bvsSjGzqV9wBqSwzk/8gpvEc/Ek
6hnfgyYCMk0MqY0CNHlq3Gtb9nSjLmZ+MmLuYhcWyfrBwFraB+8pvC8Q76pQghv0
ErN0Lwd1YFHTv2OLQO4tTHYG7KooHnS4vyul10XOC0mYJBLE8jM6Gry/7nO44Cun
LF8vyqcEf16ZKZPEQpQQlCN0pOYy5dz7El0NLojZXONRrxNn/GpVV4N4aZsIvX8P
+xo6pwETExt3vr0korpsbIUwSgWBKaXRr2/8xuQGWMhRzT3alygSV4KH3gptpT+D
IZhdExSV6tDB77jhLM0YLk/BKl67ogOt2bAF1OeH9GjEcsQvC4x7R89+8mJLkHJQ
XH3k1xc0ohcydbgX8H2baoLMRd6H9ih8a/eJG9LSzZhobgbobxB4MjWYwM7v0Tmb
VgXoirVH/lPDw6M0IilqzhElSiK22fbpmxBH44a+aNb69E5gNGeYgA/XGRYLy4dF
D4YMojPROEeZR/swtYsucaDWUsNezdiPb75dBeeLR7ZUlyEzqTqv33Mwm4tXlrew
8FR78QP9yyJvW6D/61GOHLSRt4PrBcC/1fgRDPlvRbCjLyTf+0+CR7KCq6tEc3pb
Hn4McHB/rIkRNIh+f2l8kmuz9caJOpmOjkPJlUHi2zpLUwh0NTaB5dlF2eNoO8ml
Cca3AKWylxwxo8U5Dbnjz/V6cnMaKGCXuQtivYlBiwrf/m5GfW74K4EN6tRIuPmo
OQZN+E51uEWEYI8p6qA2ihP+A4uwwzwxNNZHR4g3nU9QJJQSIggE2FlRnbjp8Nyi
zwGBL9v+HKMW34ddhYZQlNw0E2AITIuVvyM3tayEVBRLBxRQ4M3KpyPDK7DG6yvy
lBqKgD18nasOvLYnepVdknh8nS4PuikE3qwGRl350TkmwuYysHSg/T+iNEEUrWzs
yT/bseu14smV7A2/cfmMhKphWLsZXjVwGlMps0IyFBUou6c/c8UY8D7ryLDE22Hn
GAt06crr31+5X7SBOp1eXMhFH2yaUDMR/IQ/+x1H5HuPG9nn997Gv5/g9ep+XUNP
FnP8ue6WrHt2lfGq8hVP8L0nni8UPaVhrTpsIIAbxiR0FFwevfFZCJlMhFassGAt
nL1Q9+ANwPvcqlKhMM7CWn52asMW0tROKOUaZeYFNf1SPTuzaKUt4GnRYLst7By9
KtxQ7Fn8A6kUYBWSunINYaPw8Ker20YnLMEh+/IW3ILB9gq0xZykr64Iko0w5yVh
4z5wlMkWbjSo2prL+KM3RaEx8XSClMon6tushcLjI4mSaU0e2fMG77DWBxOzrBBN
gtooC01S6A+QHfH3eNHweyMzGMk3aPpp9L5HsURkorN6PzojIFUme58L0y+ZpKPs
vbBubPrRBjZKPPjp+V4yjpBsLko1Sg3sP6dvPglJwrqVifaRTteSyu+mKC53XBYu
2x4pHsmiCuqPaBuQm4+7LYhvmzUuZUFP2zOFG6OEsABvS0x5Fuo4CnTO8lUUxgWG
/xVSNf+8Vtx6kEVJhvQtCbEcy4u/j1PqtIpUeNF5jxKVnG05gfACH/ltkwzryiny
2CZ349NpDHuppUxALkw/mfIpfS0cRPIuNvcADsbqg6+r3DDKMYk0iE4mNEbGZyBw
HLjKvhFqr/DfJ/eCCD4f6QJuwht0jkyD7BTCh7l4MGtx4VctyDGHZALZ92enVDkY
A0hzI3znkJCgRaNbg5J2HoqSmzyJ2JyMF+rES5PBXISDtFT32SBI7fvi+kc76Ia/
ZvJjNGmosShDoDhRIbE4jsYZFZIPtHmPLlfsG+K0RtwMKn/7C28imwm5T/SVWtWO
n3bcYZIgaqIGYF+Tpkft/+emJBCXWXBdcGs4iGzQXfe/ZE34XolZnWaCiccJD+pG
+jpyttPjp2IiOiwf6TC5GQhYWvfCXf5znw93saaEFAtsfHig6ROQG1zTaEvuaCld
A0fEMHTRRWzoxpAr7Jd9UmrITUj1id0poEEXMaQ4eZUV+6NcbyK2oCIWnw3wD8cD
DeBQ22kCrdZR+Bztnx8vPBEAcRlMIUpJDIwoJuhnsyAD+w37y4O5jwhdryc19gYv
CVxJzHEXuvJ08rAEttGy1jcBn5/mXCRLqQm0qZ9lvQ7vTACMnpd2O/VO2UN2wTQZ
UR8DQGG5qluNBzPRtR/+fp+jB3egMgrEjaFomqP2iOVH2i6/1M+A/k3B3G29zKnt
8/Vi3jZjvDb3TPdfEuG6BokeznO4PIZoNbjl/dDCv4tmc3XlUNSjQz7Yn4h05+m4
UrZjbDP5K94bRj36l6+mKpii9h92PqE2YlGjCcGzDPibWGvZBkTRCtfTDVmYGR4A
TJDqym3F2squRL4dBeOAGAufpDUDqeCJ+dmDaB0Pg5y/QjrtxudbeovDROzA103G
ijRm2++TdKhjqMuz6zIyX35iRpJ32wVuOt79Iziiq2lcqxpGHuuoLFKqqBii2W3k
qmagrOnWqGf25JWXZlfKpjzpL6IOXWZCSK5bqHe0g0XzmGMYhagwYhqZ2b4S5R/L
+7WiVb2armx0P89EwRx+3hbgZPPeq9NVmr/ygFnRTz9uENrHy0OhcRiTvJqiVUwn
AzqjzHjnEMaqnkQRIYdaKhUi3eD81/huHlQAG100jxYlZL2z+bHtIcXgw8dCW78z
L5iir1vKslR4hTetgBz4FSFx97+MyrKt4SMZaKtWafuodd3s02T0HTF5JILZ8Fkj
N7FLY9Yr0hJo1Gg6ZfYtJmFVsPj2ybjoeneMnctetETE5LYKVM4TBprBahnF85Om
QXFlNBgdOq9asJvYwaPxAeWifW87VJRTXOANO+7OO5A/2i4TAogtlKN4y7l1lFk6
ErcxuJGv9OJj27C8xXyF5GLmDtT+mcutgbwfWySUClvRgcU1vOgAqcb9m6p0Sbme
jnakFPIF7Pc9UbFDWk3hE5djr2kvqLRwFXAVc9aKke/38rF/2DKLjt3SM50PYb7E
U5EHLn7Rna1hw1zvSeWFiiTbYh4WGV7e4cQmIS4x6Ki3jkaqDxOuerwFN25vTORJ
Z3HIqD27KetEmLmDSbPCtSMd/A0q6uXDbCL051mvg90N5NZ3a3cLEactZKHMA2ri
dpuVAcQUXowbbb31MRZLqza5XJbRnLMf8B4Fs2zV/d0LvOvnh9Q8XnCm0/sDXbAB
`pragma protect end_protected
