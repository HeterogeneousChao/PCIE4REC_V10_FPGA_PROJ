// NATIVE_TRANSCEIVER_IP.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module NATIVE_TRANSCEIVER_IP (
		input  wire [0:0]  pll_powerdown,       //       pll_powerdown.pll_powerdown
		input  wire [0:0]  tx_analogreset,      //      tx_analogreset.tx_analogreset
		input  wire [0:0]  tx_digitalreset,     //     tx_digitalreset.tx_digitalreset
		output wire [0:0]  tx_serial_data,      //      tx_serial_data.tx_serial_data
		input  wire [0:0]  ext_pll_clk,         //         ext_pll_clk.ext_pll_clk
		input  wire [0:0]  rx_analogreset,      //      rx_analogreset.rx_analogreset
		input  wire [0:0]  rx_digitalreset,     //     rx_digitalreset.rx_digitalreset
		input  wire [0:0]  rx_cdr_refclk,       //       rx_cdr_refclk.rx_cdr_refclk
		output wire [0:0]  rx_pma_clkout,       //       rx_pma_clkout.rx_pma_clkout
		input  wire [0:0]  rx_serial_data,      //      rx_serial_data.rx_serial_data
		input  wire [0:0]  rx_set_locktodata,   //   rx_set_locktodata.rx_set_locktodata
		input  wire [0:0]  rx_set_locktoref,    //    rx_set_locktoref.rx_set_locktoref
		output wire [0:0]  rx_is_lockedtoref,   //   rx_is_lockedtoref.rx_is_lockedtoref
		output wire [0:0]  rx_is_lockedtodata,  //  rx_is_lockedtodata.rx_is_lockedtodata
		input  wire [43:0] tx_parallel_data,    //    tx_parallel_data.tx_parallel_data
		output wire [63:0] rx_parallel_data,    //    rx_parallel_data.rx_parallel_data
		input  wire [0:0]  tx_std_coreclkin,    //    tx_std_coreclkin.tx_std_coreclkin
		input  wire [0:0]  rx_std_coreclkin,    //    rx_std_coreclkin.rx_std_coreclkin
		output wire [0:0]  tx_std_clkout,       //       tx_std_clkout.tx_std_clkout
		output wire [0:0]  rx_std_clkout,       //       rx_std_clkout.rx_std_clkout
		output wire [0:0]  tx_std_pcfifo_full,  //  tx_std_pcfifo_full.tx_std_pcfifo_full
		output wire [0:0]  tx_std_pcfifo_empty, // tx_std_pcfifo_empty.tx_std_pcfifo_empty
		output wire [0:0]  rx_std_pcfifo_full,  //  rx_std_pcfifo_full.rx_std_pcfifo_full
		output wire [0:0]  rx_std_pcfifo_empty, // rx_std_pcfifo_empty.rx_std_pcfifo_empty
		output wire [0:0]  tx_cal_busy,         //         tx_cal_busy.tx_cal_busy
		output wire [0:0]  rx_cal_busy,         //         rx_cal_busy.rx_cal_busy
		input  wire [69:0] reconfig_to_xcvr,    //    reconfig_to_xcvr.reconfig_to_xcvr
		output wire [45:0] reconfig_from_xcvr   //  reconfig_from_xcvr.reconfig_from_xcvr
	);

	altera_xcvr_native_av #(
		.tx_enable                       (1),
		.rx_enable                       (1),
		.enable_std                      (1),
		.data_path_select                ("standard"),
		.channels                        (1),
		.bonded_mode                     ("non_bonded"),
		.data_rate                       ("2000 Mbps"),
		.pma_width                       (16),
		.tx_pma_clk_div                  (1),
		.pll_reconfig_enable             (1),
		.pll_external_enable             (1),
		.pll_data_rate                   ("2000 Mbps"),
		.pll_type                        ("CMU"),
		.pma_bonding_mode                ("x1"),
		.plls                            (1),
		.pll_select                      (0),
		.pll_refclk_cnt                  (1),
		.pll_refclk_select               ("0"),
		.pll_refclk_freq                 ("125.0 MHz"),
		.pll_feedback_path               ("internal"),
		.cdr_reconfig_enable             (1),
		.cdr_refclk_cnt                  (1),
		.cdr_refclk_select               (0),
		.cdr_refclk_freq                 ("100.0 MHz"),
		.rx_ppm_detect_threshold         ("500"),
		.rx_clkslip_enable               (0),
		.std_protocol_hint               ("basic"),
		.std_pcs_pma_width               (16),
		.std_low_latency_bypass_enable   (0),
		.std_tx_pcfifo_mode              ("low_latency"),
		.std_rx_pcfifo_mode              ("low_latency"),
		.std_rx_byte_order_enable        (0),
		.std_rx_byte_order_mode          ("manual"),
		.std_rx_byte_order_width         (8),
		.std_rx_byte_order_symbol_count  (1),
		.std_rx_byte_order_pattern       ("0"),
		.std_rx_byte_order_pad           ("0"),
		.std_tx_byte_ser_enable          (0),
		.std_rx_byte_deser_enable        (0),
		.std_tx_8b10b_enable             (0),
		.std_tx_8b10b_disp_ctrl_enable   (0),
		.std_rx_8b10b_enable             (0),
		.std_rx_rmfifo_enable            (0),
		.std_rx_rmfifo_pattern_p         ("00000"),
		.std_rx_rmfifo_pattern_n         ("00000"),
		.std_tx_bitslip_enable           (0),
		.std_rx_word_aligner_mode        ("bit_slip"),
		.std_rx_word_aligner_pattern_len (7),
		.std_rx_word_aligner_pattern     ("0000000000"),
		.std_rx_word_aligner_rknumber    (3),
		.std_rx_word_aligner_renumber    (3),
		.std_rx_word_aligner_rgnumber    (3),
		.std_rx_run_length_val           (31),
		.std_tx_bitrev_enable            (0),
		.std_rx_bitrev_enable            (0),
		.std_tx_byterev_enable           (0),
		.std_rx_byterev_enable           (0),
		.std_tx_polinv_enable            (0),
		.std_rx_polinv_enable            (0)
	) native_transceiver_ip_inst (
		.pll_powerdown             (pll_powerdown),                                                                        //       pll_powerdown.pll_powerdown
		.tx_analogreset            (tx_analogreset),                                                                       //      tx_analogreset.tx_analogreset
		.tx_digitalreset           (tx_digitalreset),                                                                      //     tx_digitalreset.tx_digitalreset
		.tx_serial_data            (tx_serial_data),                                                                       //      tx_serial_data.tx_serial_data
		.ext_pll_clk               (ext_pll_clk),                                                                          //         ext_pll_clk.ext_pll_clk
		.rx_analogreset            (rx_analogreset),                                                                       //      rx_analogreset.rx_analogreset
		.rx_digitalreset           (rx_digitalreset),                                                                      //     rx_digitalreset.rx_digitalreset
		.rx_cdr_refclk             (rx_cdr_refclk),                                                                        //       rx_cdr_refclk.rx_cdr_refclk
		.rx_pma_clkout             (rx_pma_clkout),                                                                        //       rx_pma_clkout.rx_pma_clkout
		.rx_serial_data            (rx_serial_data),                                                                       //      rx_serial_data.rx_serial_data
		.rx_set_locktodata         (rx_set_locktodata),                                                                    //   rx_set_locktodata.rx_set_locktodata
		.rx_set_locktoref          (rx_set_locktoref),                                                                     //    rx_set_locktoref.rx_set_locktoref
		.rx_is_lockedtoref         (rx_is_lockedtoref),                                                                    //   rx_is_lockedtoref.rx_is_lockedtoref
		.rx_is_lockedtodata        (rx_is_lockedtodata),                                                                   //  rx_is_lockedtodata.rx_is_lockedtodata
		.tx_parallel_data          (tx_parallel_data),                                                                     //    tx_parallel_data.tx_parallel_data
		.rx_parallel_data          (rx_parallel_data),                                                                     //    rx_parallel_data.rx_parallel_data
		.tx_std_coreclkin          (tx_std_coreclkin),                                                                     //    tx_std_coreclkin.tx_std_coreclkin
		.rx_std_coreclkin          (rx_std_coreclkin),                                                                     //    rx_std_coreclkin.rx_std_coreclkin
		.tx_std_clkout             (tx_std_clkout),                                                                        //       tx_std_clkout.tx_std_clkout
		.rx_std_clkout             (rx_std_clkout),                                                                        //       rx_std_clkout.rx_std_clkout
		.tx_std_pcfifo_full        (tx_std_pcfifo_full),                                                                   //  tx_std_pcfifo_full.tx_std_pcfifo_full
		.tx_std_pcfifo_empty       (tx_std_pcfifo_empty),                                                                  // tx_std_pcfifo_empty.tx_std_pcfifo_empty
		.rx_std_pcfifo_full        (rx_std_pcfifo_full),                                                                   //  rx_std_pcfifo_full.rx_std_pcfifo_full
		.rx_std_pcfifo_empty       (rx_std_pcfifo_empty),                                                                  // rx_std_pcfifo_empty.rx_std_pcfifo_empty
		.tx_cal_busy               (tx_cal_busy),                                                                          //         tx_cal_busy.tx_cal_busy
		.rx_cal_busy               (rx_cal_busy),                                                                          //         rx_cal_busy.rx_cal_busy
		.reconfig_to_xcvr          (reconfig_to_xcvr),                                                                     //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (reconfig_from_xcvr),                                                                   //  reconfig_from_xcvr.reconfig_from_xcvr
		.tx_pll_refclk             (1'b0),                                                                                 //         (terminated)
		.tx_pma_clkout             (),                                                                                     //         (terminated)
		.tx_pma_parallel_data      (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.pll_locked                (),                                                                                     //         (terminated)
		.rx_pma_parallel_data      (),                                                                                     //         (terminated)
		.rx_clkslip                (1'b0),                                                                                 //         (terminated)
		.rx_clklow                 (),                                                                                     //         (terminated)
		.rx_fref                   (),                                                                                     //         (terminated)
		.rx_seriallpbken           (1'b0),                                                                                 //         (terminated)
		.rx_signaldetect           (),                                                                                     //         (terminated)
		.rx_std_prbs_done          (),                                                                                     //         (terminated)
		.rx_std_prbs_err           (),                                                                                     //         (terminated)
		.rx_std_byteorder_ena      (1'b0),                                                                                 //         (terminated)
		.rx_std_byteorder_flag     (),                                                                                     //         (terminated)
		.rx_std_rmfifo_full        (),                                                                                     //         (terminated)
		.rx_std_rmfifo_empty       (),                                                                                     //         (terminated)
		.rx_std_wa_patternalign    (1'b0),                                                                                 //         (terminated)
		.rx_std_wa_a1a2size        (1'b0),                                                                                 //         (terminated)
		.tx_std_bitslipboundarysel (5'b00000),                                                                             //         (terminated)
		.rx_std_bitslipboundarysel (),                                                                                     //         (terminated)
		.rx_std_bitslip            (1'b0),                                                                                 //         (terminated)
		.rx_std_runlength_err      (),                                                                                     //         (terminated)
		.rx_std_bitrev_ena         (1'b0),                                                                                 //         (terminated)
		.rx_std_byterev_ena        (1'b0),                                                                                 //         (terminated)
		.tx_std_polinv             (1'b0),                                                                                 //         (terminated)
		.rx_std_polinv             (1'b0),                                                                                 //         (terminated)
		.tx_std_elecidle           (1'b0),                                                                                 //         (terminated)
		.rx_std_signaldetect       ()                                                                                      //         (terminated)
	);

endmodule
