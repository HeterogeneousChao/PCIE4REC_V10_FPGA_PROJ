// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:19 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E8gF3vXoRqCA8bE8gPWEkLZST9n+iOLFtQRb/pyqtkCNCmFpiq+q2Q1W/O12gBTb
uuC7T67saCT1Z/tKsAWj+WIF/DXPDiHZElzcefCmYhJUwwz2caZRPo7K3SItJ/Yk
sBmWnzSV3IJ6tjsNwH6olE/W131ugTMgE5hMyYRaiic=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22624)
9cMb9M2oDYI9YCmqS7cnkma1PgV4b0FYx7clcreWt/yLspreJ76b+RSVULGF+ojQ
K11Vn0AFP00ugX2Y/rCBnXayH0LrrUi1uAarqCMLYOAaY7rQ0uV4Sh5nlllNRNYS
ooiJfYJ5bDN9iDkK8Wrdgl/eTmwr+EiBXNZwgmSG9zEQgrrWFjt7RzScUrycPWKx
MXQRPYn4EWD/V1GfGqFuw9DR4fyi2Rw5DkCW/P2eVK90K/KPnu01oDcSlvQvhVB2
vHNAWLDbEbylSBUpfJGVT6M90YMFm7NUtxdYi/b9qTlMtJ2XzWA9O+0F16oF7yTp
qZuoVD/PxXBU+0AUS4vg4vRxYHjzZsm5ZTKsNAvM16rI75AZSj3iok5gymmYAFcn
TlsGBgcXl/ZP5RL7KT7YkNilU4uKQUH8dezw8I2L0th6yjxvRSTbwDFemjMHfZbl
W1cynTJmrhpva7Bti9UySCrM+Yr4UIi9FZ0cud5efLnzg+lw7gVYaYJJu6sou2qr
fmjMRjNv4sfXdAizNUXftUFiZ8xE30y3MVcIhzhB+Tn5atZ1WjwufIM97+rKQeyP
W5OOJS5SbP18Y9B8H+Z+cb3um1MUCUAH2Z5LMP8qG5jCMrl3Uvg/liqnclmyiC5M
8WWXjCJRem8V7laVdUCICUmcELOtRK50i6YFJzTvjAVQp5Ps5uHHBXoIjkpRlauK
VSUOknSGK7JVoAjFxl0djECEyqZLquY971kcoDeRlv7JJhI6jhpm7kzdQRqPUUG/
EOtTSiTfXB8BgOES3N+uQpEW5Zm56EqpLW939aubk68dlP9BMpgDJRfn58R7tSto
YWPykxjZ14q8q36HXJxTKHm1m6j/eJtXUiN6whbi8iKA3nlviwwXFt+4vfiImwfF
c3iqHRXdJoDX9XvIHRhlbQmZuj8ojLPRRuRzXKfgMp5CvgNR6Xa+9s9JHwx2zAHY
pM4/eNqAsZRd//JrJgEOX4z4y2C7CaPHtVhebl1RUuK1ewXS1DndyYovvnrTm5j/
LRdJTS+qflFgG0cdQDds8eVr7nTmZH8XTGhB6om9xj76sUfabXq+LZHLYT+c13SE
6c+lAlWZGtcBdMcZaeSk7zl4SnS/juDLN8xlaN6hevNnoKAOJlCp3eAhcxFteMue
Xm+HyiDYqEC/eLuw3kgSO/Vs59jbDz7Y4UXawOIi02LTlCDZyip8SZVjHXIA5M0U
r27J8xHxejURQ4XdZurMPfSIum17R62roncD/VcIAPR9x1jAYs2uKI+jTOJDSZhW
L2UPFMglvUMswgy5golVoEPGZajnOdOVbjJa656bzbJcRl5eCUUoaWWtY3Kh6cUe
6tYJrxctAgLYZBlfhHWtAVofbBFxrJy7o3hKCfCcScQ98rpNhE4jvE5HjGSL17Ip
CCgdBl2sgBd84Yx2NQwSqo0wacw6VqorfWC0/XvTxPnjYASEV7SRcNFOqFryPvYu
T8U606jNdPM2b7p02Qlzf7CkJv5Mz61q89LOXWC6yqYCTgyEEcQtvDdU9nPFlsMq
bMnOmJMjtP4GXZiyF3btFgssb7HT/TvrcfPwbXbU+oR+JzU1ygqoPmYnhWZaSCEZ
RTRsjf6DZVkkngmTGBt8S6vdP1VvAmNM0bfquXg6WFMX6NhIvDhm1Q6S0bvD28RJ
4OA2B2zUKbusOVL7j6kuSZvIMtxRR6UGLaU86cqfXSssxFQhM8Wt5yAFRP4ggNPc
ucYEYxCoZuQ0iFNVbm57jBlTi6L50s4zPI4EIuao1ipB7BS2chyiUXE7MMB8TUV5
u51HCYHfGxaL5ec6sqTqgzaY2A9pSlJY9DKb12NwSinwac/qkq4h7MOtDzV7nDRy
8VzeMaoTURyTHPrkcSD3bO/+kbBFs5q9dY3T6hj7DByxW4BIMqnUHwxLP80mzkJO
NOV+VolKO50KVaZ9aUM9XVXGRD62hydzmj82IXfQ0lQT9MO3o+cC6J3UkyiGa9W0
O2DFpJCdD2biac9qZhxbJ2gRjD9q8dRIyJed76sW1T8DNBcutLsqdRSM65UlCA8+
GxRXrwUrLkvqNEj/6QRr4xUeAUFWlltoud//sr5AouzgIpjnMAU+1Cg8haoaex3K
zcyQF7XYA1y/0K02OvowM3HAunMZAVVxTt/SPzHjjPVZU3AfocJCrmrXGABFY0Nm
UnOW+HedaPACmUPZnal4ADxd69yLPAmx2cwmf2njD4+cbLnSA4jAKmiFJm3NCfZ8
zRL3td8msxZlEOqyeqjnat7vr2Gfnren1LcwvFuHkTb+4wimVMrD4KwAcjVNuUjd
DWovV26NXQqJS35OKlbQrA07ZO8NHvjoh7s1xT4SIl/g+X/OGqfQgPc/er34+9zs
K0Nlxn/jL3UIbRWAr42175P9Lp4afwUK0Tljg4x5hq9hbXfWdLo4xv66BY99GJSc
518FANvPp5IBVAin4YlUi7+VRfSOmGrA0Mvu6q2t8ClvxOB93zBI4Hi+tiG5I8Rf
VmVx531YjCyJoHzkGsvez1S4m/5Uqg2/frZlzCCZqrl2b9EnTGVJgE5sooMFBXbh
Ph2yPWLX5uXV/G6vUKWtzZmMkRcPDCx7qyjmD5HWTqQ3ZG8odA4kYPwkxfSL0Gp8
et1Q40dHPLO1QaVIlIvAZF+ApxbaDM8ZovfOn4AUwckV2kSNqhxpdhdruDU53oaD
pxnrEnOHuY+SA8NiFjvq1SGSppZP6w91/y9/GxzYV+rpvCWxKVXuewhZ1GXwXu2n
LVA/JdQqis17Vw+/Rhr/LcUN4Sk9dmETBONuy6UPsFl5G+UrQLbH01qbFjvhDdFa
r5OTCc7U88R2ZVyFPfwkekHF1lD7hopN+dihifjsxlW8tJGNlMhYeQG3riQJRkNJ
NddZ8bPBe8XsMkbrQtlhN59i4MIwEC1M8e1PqGZKIF3iYGU7snuOCnlayVRhLzwE
I09Xp3KS6sqUEXSOoM2r8wTwTCAHgdMeYBc2BekwhEHN3ViW/uKt30bdNqKhVHej
nO1JznGUdC1LxAfGmzoruEwyJAYbED9SMOdUyJaQyKYjHzWsfrNr6ivRRL5LbK+f
sNZ9OcoTGvVGAmNPU3JaUmlzUsVRPb3Ad+RZPT+3NfylMrYYd/eICAIQLa3DJ4UT
v4FQXU4c3lbskIrRhmW3E1bn1/yzFRHZEGlm5U1BLk9JRvFjUkxuNgBiMGF1ROwG
p/QR2UY5GRA/YefAb2E9PPt7igclGCv/Hj1DnXmbV96DEDflaDy0hPGNJ7CQX1Ih
When1ypMtePzVwAdcODXtfbS0LTh/WxpTP3ZwQP5d6HjGy4KkIO6XmCHxqBfhFSn
Cm0ClL1eTfVATMgBm8WyvTrMr4LK0Eov8wYGZk1GFXFH9yTpWS6JxBQVYnN7Owzd
ESAhny8gtaEkicYTA9F5J5lTIrmXpcdHY6OEMyBs1LBQSO0eyXQsGwMhE3E5Yzj1
em0XUEXKF3GTEtD1t5CyZOG0xsUhfeN4olT5EiqU8kChtGbl2Jc/PCpNgfozcb6u
PQZ6XZZ5IucPSzmBnwdegPH7uHzIb/B6XuNFQtadhpwMRA4bpVT9XVeGsQ/hqsQc
RO3PcWQhYnj+ooYhDDRzJYS6jgGnW6flY6q/HJXxJnPej5iTqjDjeTO83Isdvst2
U5VfZCVuNDHb4lShk6DN4ITLvfRLkHkIKSTp6oCRSxh1ex49UYLDtyT6EwP7ZYS6
wNQolTy7ci5+lIx6WRpIBJ7ngUvU957TSyL0PUlULx/RJdy0hAHwVPJfvsutBj4V
Vhv3Hdazl1znHA+w2bAOtniobkb1I4GVWcdcUWruyCymvW2MiGRuYKYiLRmdPGwQ
zkg2VmUzs3cD8RfdokBzJ2j3NyOHPr9ZFBfevgFo/mZpLkyGs5XmiN+rDQ5MQM1X
XiojhMcxti5+Q0DsoZZie+TkqYuhTKmYV0qt0ZuuTX9d2JlVB6rO46Qj3KU1SzJN
J1JREdmcVD3Q+KLZ3tXpkGUSE2TsmQqNSQ7+MTAfqc1CZrUfy38sfrHHYKHTSa8j
VcNBrjYvI4EzDPpExzzsVQ6MaAbwy3/WQeKiI/6GvMjHq5T7GmzM0UAeXAeH9lu/
LGNAXdg12s1sMdD7mxF+f+JYz5EAWO1Mb+drHWZkHSEZ2FLpm6e7g0LAr4OVoXAa
/8Zod+ScGDJlKZdG4c+y/nvtGU23mcMHzTxEZQINLr42sFJjHPLl1Ogo/DGKInCy
z6ly0Rt/je6ctkpCH408l2I4OTPM+Z+XgqDEsGWeDOvB5Pu7ziIy4PhnaQHOEpqd
VeShIwBBaRbclVdi6wEWGCmQK1na1gI0lzhGJ4Gb3ihBiW8M/ueR12e3pUh3JTqy
/PF5tEzqy70YZujbOG08Ujc81uvdnXZJo9m683yAXltU6hlo4M2lDAQPdUDUx0S7
xX/JxSgTQknW59iExVLHUMTMQiQP7BefgxZXQZ5HcwlOPaGGPRNKo9vvh2g0r8zN
Cap1nD4DfuxRWQALR5Z4ZC1epoSXOKyN7eKO+uFKP9WOu1/4wYI1hgn38/3cB1sb
RpaXP/7VTz0J0bA7ljrf6QS17Mv/ROcwtxcqgh3HtxmS8ZviCE62iJlqR8t/Jm9H
Pj2rlXUCh7VZCEPzx/GhSbdkIv9OnKu3LhK/ddsJZap0d0QlYDVHIUjeGGCMPBkM
xVPXhmGcIisaRfkApWVCCK7S879OfbnDDvA868ouQATCQRIpnxTzow7wXFsUjTBB
qPwpDMoKHRv9JsSMJcFNZ4E9gFUoHnYHqtJW5OR0U9/G4IIje5MAaRGfqaUIS7yC
xlQzDw4CwKSlItiLyI8oLRGbnI2W4o5Dc+2eJG8al9dwE0znKmpcoXWEIyzCdp45
fXJ7x6/zl207D848JsZd0yZz68m/+JzKAtZr2PvLKVAPWS53LEuel+3DCJ6t8vv3
zEIKZzd+kFv2hMwqcOP1y/DX7Yza6FUna62nZY/8kkH6zrZ+6rrqvBLt/DImQSL2
zgqsQxZrc93qwaj4MOPWqxNZMLZsUsVb8Fbb1IVtY3bAxJv8l7E7eOv/ZrApCfxV
b69JJL9sQKRPHPHUtsv9PlxkFpUgM0YD4cgEr64IKExVVqj9aH6BAOUwJKharzv/
FAyveBAn3bVf7UROwd4YvANgL+vKVfRXClATC8JQs9MRCJyAU2Opotk2DtIpi/iC
uMTkQrz0nfAOlz0nNPuj6Oi0jpLNTql/m7s7yCS3VbEwtYue2mDFmZ46wDdC2kZf
ItkQcXZtDaEVeaR7khAsJVBhXW3HoMNWYb3+0h5zQcbw80+6ufcxdI+Zwg4QrJVK
eradjB1xQjk8sqSln/yMZPBLQrsIqrrsdTRYm6eBHH83kT10cdj0O6ZpQfKCmDVp
26bS0JC0djFk5KuCYh5d1geTcWg6o6yKNqMpSmw6eREM+XvsTnpiduZaVMQvRW7M
vQ/n4d30OYpLz6trSFjYlCN74kOTuQ/76xpqpwPllmYiWFjfYj5QXcLj66a+GRRt
2FlXysIKmpdukLqg3E7Gr/7mfE5KhuugcJy7tdh0U75R1vuKs9/c5p18cvt/K/Ap
CwY0NFsxmT9Mj9JvG+IFuonaHzdGVR9X9uafKxkBPHOWpc66og6H5pmb1A8DRSzz
0/LxLZhB/IoYdu2kCrY6VATgvtLi9ze88jc0hiDDOlBCssNG3/ZQ9Wgv+9hveiH8
Zq5UqyKrYy3yxGaTJdH7u2+MVHYfd+skvvnop5JZ3Ml/o1TloVYXWPsrZ1aC7x7H
sc1FGhYku55hPYnr79h/2lWnqaHg54dlfMInHf7ZpYshA/cTr0lqntZszEy2hFBS
y+uY3jUkimt1+QadIeVIxEy6H6oyCQ/MSJ+wfs0rDegvO1I2A/KJZNu4khZas2no
wGzotBzlA0FB7gwuEqXY+Z8RkeJOhd/zjnIZsUjc4gF54RYUo2MY8pXanbqWnOPh
1s59dy2qZA2tw5T3PvyUVyhHNn8EIGUj+Kph/tApasAxULDCTxNAuKuZOiiv/y3J
RafrzXHrEsB6pYEsSQfSYjPSnefwRPMiooJwKX+VgHrJBTaf+YGWCTFN7wjB/1r+
zfNgaWWSvXfkF2n7FscGbAF5u686J6yuU6EntvhkOrHZ1xKTiGuVTJW05jUdatZV
/fKy3xhKUS394WK0jgOjjqav2naRMYieoOjaON5C1FQ8SYGXpQmPPo6OORZrK7n6
YXnm+CRQ89KCraqPiFbg72oUVd2AclQTA7pSmRPsyB6q1ZG2QjJfb61rOwIxZZhN
Zq8Bb9r4xF4TQoODLl2NjlOfEouyqNrkRXK2fa/TO9zI/8y9ul5ql0wuxXrU+t++
j1twxAPGjFZ87q6kVvW25XQwAD+8sBBOoO9m66RO8e77kEswR23P41vnWChgz/tr
Ycw5n1nvCne8UsPhP43jxqlNOBBN1YU27ivWieTffDa5RW5W6jHRZ+Pw+J5w3v5O
K/Eh8LREDete+D01XL+Yl8Fwf0EoT7pLSPOOqbGkgWJIrfmpBuDh3XbtU7zUYp9B
d+Fifx5hUIQKFZbED7H6uyoe+Gqob85OQJPeVDxDRKwg7Bj8ghRFeo+pX48aJc9b
410qFN/yGx7j9j9EdXNlpBtoJfIprtLqpMP4SDjZE7pfShOzVfce2Q8iZBxtPrNt
bnMIF3RBki2cJJDBckmHiGWHrBbfL08FK7km3UF58kyF4NDcJ2eJYzrKQtBI+ipu
anNbyMZr4fsScYgObf3WiTx98PgpjHpqRCJTHfudCaE2R9YIujBEjZjRHxKEQ6Ha
zL5mH7VtJQIEty6bSsnbP9iRf3UoefvyisG4bKX0TLHAKc9uwHtsdI0TVbcOhh9F
mzvVTzPeh7Fgj69sWYF+UZIE7oCImzi8Qc8rjufzEpPSkZyiAPJ64nQ1Z4uikhkY
AtIDxnOCJMYaSmE01ydEzXa8w0dTvtYE4m3b43ICQ5bGhczio0pq1TqPEOXpnQBG
rl/Y9HID/ufaeqeRWL5QoYeNpIl2vZVA/9QBQPLvDq/NSV+B3REGXX36sbKYfYUH
DKykVZy+1iP1K72qxdY2ysBkq1nBn02djb8FGz0yA3IlAaNwHIN2f7s/ek9r1rdB
p12MJMlWQpyg3W7m7+YwF9savij7DRCZQnN3DbSoqJrWtycMhfvaxJOmlL9n7cCV
gnvoWwrMpbOTl5gRc3zB5nGuihEhDoBQnQ9hA4a6eAyLDKhzdACty5qRCAgSlUVL
JS5hy9VaozBwf9WEa1SoUYvuGYbF5Nap1KvuDmesWVC69fH3fm88YrghDwLJac1g
mEAY/oIB33vvhos2nQAll0ZE1haevsCyaBqU2QIv0ZXzr+E8BKVQTKugnP3ahGES
8btvBmcGPHI7NSbg78VPutaAU+2nSTSOrQ8nlNm5dfBavolPAPitD1fPbF8h6V3J
4OETJvtoN7rSmAt1CuHgnsUEBSy4CSh18C51xL+2zB7Drk4vMqcyLxHKZ5rcq/9k
YQ1c3dYLiIlk+/kKydJm27gnTTHQlesuoHWpYTZiJp0Wp+aV6vfG3/N87tKWB+Mi
PRgksufoKYB3Wia7T61QKVYZ7/zrLE7+40DxirVNF+TEjzA9i0pP4Ot42xqXlxXk
4qrjxMZtSepxsSS7KSBvvalmNxeHJpx0G1HkF/eKMT+4X49FIPPFB3kzqWANcv4Y
AYVcYafzok+mYMH60Sd5lSANKxf34brNjXbjYZ+qJrykYii+Wd2QkYqAY+ZuZlQE
UipRg3x2sWZLDYNW2oyJYRkOll8kD+mt3tZurFvnAXTSwhjKevE7Is+2v59oBtCJ
7Dkaqe+mUst7QAz4I+9a1mrvU6YnnHfKRhMow0Snk726YktKy5TJ81fDp1Fk62d+
oRWXXj8KtA08uz/HQ7vWrEvFq6rq8u5s11ft4fKFHvvGF+uyLqFSW5KhocYqKPNm
dY/Ir5vuDfF2JnBO1K/xP12h5HGGS6yBFdNnX1pURH0k0M2YV+26L9JX+9XZDtfk
IuK4OiU7CZzXb9E+iLOnAa+trJ27CwfcYW4bESqR07k9dtpPgPQEjt0kFJwFJYYr
TLyEYT9mbgukpyRXnIMBCd9kU6w54Wnwv2Zw1X1PgGkUQL2Paaz4MhTWt7QujCfD
bUq+FDbkA/Dvj8TSjC3KcB4X/8etXRylQrnu7arZBljf+ft5QMgmrqDgaIW8LGE4
fqy7ZsS2po6OKY0TPH0iYBIdl8hdENXdHp3xEJSUgcx0om/pE2MeR3iFQRO3karZ
pY7TniXOtP1oSYBt1b0zBlMJUsyih2Ahsft2SQtAV8D37DKQq6oHQDzCv4/+2tJl
P4ZfBldfP1vGDe+xoUvnk4ceZZ1mEOgBYvlV6gO3LxsPs4rIUn7eahZzi5eUOsRl
yOoAGwl7sVZzYSbmBy57OKApaQL3RM0oXn2j5xg+nC4zOQP+fvL05ySe8msO8ryP
wt+VwPw5skAGP9qcERbEIVOsuOp2jiIkdzR1YhDEcTB/RlzSERvOCICq1l+dbnrw
ZdKynkc1h8thH0jr0xK2mQwywPGL6wvFzVRIAA3Wp7oOqVEOjNwERLcW9Y8pHSds
rgJndhqg93rn0OiI8tSKzksjK8t9eQWq9hiMO6gBF7d/tj14A57jarxEwyTpF2nQ
v/bxALs+zNcwQjU7z+eAoqpex0DK3GkbnhGkdSgvvDY5CTpvLxuX5ZmzjBOEevUH
NMCSIGEfZH2sgtHr8xuDpJ2htCe8kpFWfPwcOVLnpydcHY+2lPQ2GepDVc/EoN/B
8YmHziXOfa1vEGJniSFVStlbE9G4UYqzRVFb67nuQ0l39cvNWD0+/oC7L2CB/ICE
Cg0Mh/Oi/Tgem8mdIaQ/gn9vaShSPhVLtQ4bAgoD7QnSrtkG/vLJXD6FeiVgE1V2
VeKfDescJVjZwKzWZTkhLS+CAuzK0v2kLITiIGIVLYBLRY04aj7nS2rx9TPaUhSR
BwDW9F1WmMITzOQzyY11Et456k/F24nAFlRV4+XEpD5Jyey7S7hHHmfGF1rzEvHz
e5QxoFF+J1Jd34mnxEBFIb+owH5WJXh+OYbaOsTd5jHz6Xe2fSlW3IQmzqhJG3XU
g931yoLQLImrHnB3I13kjj3wEH9kH3vbMuS+Zvl+JPCMalahm3Zyn7wq5BXYdDb0
K4c4EmpXEAcXw3+kB3GO+j+aXawkjmS2VV/0R2FQsuGpSEtU/KBqEXXsX7RAirxl
7gInGT0DkvVaI+9Vd6TRU2Y33548UhnFa2PtSBR4MWkAG0ZPu/cNe65crcntH7dF
ho4tOxtZ/Kto3qxUbpTX98Ej63R+yj5/OqXN5qSVNJ8OUQfswHJWQUovnNKmJBEY
T1trZjw3/wxfvLfhtyvMKzzEclzginQ6x/Zp/CAbRyTxelUWGy9zfdj3ibW/6oJD
W03E3/6I+YYQ/j+3Yrmw/npPnUrruo02xihLtd7WQGwbZa+DMlSPBXr2UJDzv9So
lFsovSoxgVM5I+lHwgMRHmG19T0DG2imdTbZTG00Kkl26Hegn9KyHEfn5yHxLfgl
O0OaEqVaUpMHsMmCKE3js41YscyPsmyh+GfsyKedQKBvlk+jWostcwyxiuXx3dAV
f1YK2PD4rnDCtsvKk/BuPv2lP9QV4wVYs+9CbdHWFkU/YLWdeHNaoATk8hIQ7TDc
ybYra48vYzTqRkLkBUpi0pVqFlcEkkIRTGhvA6ZAHgayoLWySTDgI91S2DRH6tzb
aqCAxzYQ4t8R/nplnRpjneAKObbgcPJMvDyDiD+x+2uKIDVrO3Fy3h0Ius0z1XvL
kSpQSsh7OKQvnWCTFbHYosoYRWHMWEUwRpHUMfGsXk+nLj+qJhG/5yCpYld5fGek
yeWt9rovDuB36k0eJpUXiyvYo6ej7YjBu6cAuOLgboSW0naBks59GnfdE/Z/JzSn
mwda2eRNXg1oW9Rp2YVi3GqIk8iPFp/4j2SS1xKo2EYRkWcytaXDbSiIVNBMs0lD
+obXLqrxdusybA/+kGhovw/GEvyveHvle+W8tjyTfyO9DmU8pXCDsTQ0234zrQDK
WH2YZfmVVCwQus8RkrxwFZ7q2ENFecCHmD3eEoWPx7/WKMLcK6+g22L/1wc4VIjC
FlwujoLTB7tZhjyRJCUi/+Kz/G6m929JyE4vJ8tzOy+eGG4GsDfRatNRyy7no2U+
LVVjuOjpW6Q/15hOSx9JVuLSjHHplWmCTTY9toAyLKmG0f6TwcdMoXdOlExNy3Di
QWDNWikDnRhhlH/Cy0FahavJ3vgnq4gQBV26t93CaxHnDJCDmUlum5/4IEBTaFjF
ftoxTKschlR5W7/XQUCTllRtj59BRBD04YD7PruXvvDaz3eHwwSTyKoQbVu8pzK4
apAsn8+i9QsiMVRSbo9ropXYX1ZJ3SD3bIk1vy83SgMZwn8ehhDUhbE3kwwLbS3A
BNPYIePUbTE79U7p0R1nZAavxf4ZEgFGBwpFUydXmNt2ssqBSeNWylvixI2JFCwG
wE4/wg/e4ykrQD8ZL+XCsL6PrihoaJTMYdFK/MfQocbKay0rYxzmsYD1VSUADnoN
pkp3rnVm8v7pNp9evVsdwcOu4bshCnwmAOEN3ZPaHXbhv3lwc5VGJoEQXQodulXk
ejs3gtN2BEwKxn8k81IqzmVIMj08FG38qgGD5VTN4st8+RJAA+jz6juD09soR2jq
BImT1y3m10Srp7MHsmPwsAUN2iLUcgSiUEDWgJ0UHgGxhVu1D1Xmq/k/lgusuvO+
0igbXl6kR1n6lWqD7sBiMf3q7TJvMgfB+CeWq7u3AnJe0czCf/ruIl9L0ZmKjb/8
8ySf5gAh2yLxOITavkTPqW2mQvZ4z2qu+jfFINYe4kD+WEsWWGWDBlTD6PHYyyvI
GJ1SWAL+Pfx9B93he5E78yx9hMGznq7KFojq7wPIaVRgfZ4f0LPUrlUVIy3Jt/J7
qfTs7QO8Dt4pVwwjc5CQgwKlILBLTSSt65CyaAL7b9IZhF84o8iRXBbg13B1Hhkk
4peIFe5slhZP9e6G3ZkE/qOF6pkxbVzt9mum+JJUOTGnnsUabf59KiIEupJI1P11
0ZXk/k1R9YrwW5+EtaAsg8ACqi63EevVO11VH3cIHKzOustCm/UX43R583E5EzJM
o3jHumjiaAq7aysb837Qc7yHHQrZftDv+rBs2rwDDibkPNb2vq+bGh7URtgZqcUw
ip6V0H5/S1ZGIQIdeV/dxU2q/Hd9P+0UwzsUDeodDUsm2ADahzJey5hjjrt9zQrj
oe4Ag0Z/YsicWE2n7b5j8OruGfGgb5ZGXpBsub7EIoKoAw8uzYItXxWYS6vH/qty
+nDI5OXwdL1Y50KUU1S/6CSV9FirpCcpW/ZjOoR13slJxcqZsnUVzFuohrJmfJcv
l8pVls2k+xcoIm0AuiWvjvcdbXE2G8hd1sGA7fAbhObV6hGBTskrydG+/ph/GK5m
0aEWLVXKoZFfQMvbfB8WjrO8k2aUsDP4hAaLyDb24le+ZndaMzkx4PJcAUNeYiUp
7AFfBGlCN1+b4IOfqIhIj8JDXlsgQ2DfgX9UIYGc4nsbj498+JnOk+bojzOaMVwk
TFaEqE/RI7ypPjFX1EFI8/TMCz3WcjFjwTYXJphKQay6+9IYITk6ilBqmQ20VPML
NEVoNYaKrYjbfvi+0mf19WjyL3jz7Vt0gVggUodnNWKpzOUWx+HcfCu+TG5Ag4ej
a+ym/IHODDM2nJ39VdS/YQ9a6mhvu5FUfA1h6GTquMToyOIHc25dYOyKibUY6KR0
d1MKI7zgAUWuvKHxsyAdRSWUlrl/ZiryHNmbtP+V81BQ3ilfdmY7+sJeZryAVM99
DqOmE2XNSN2KrQVIQbueMwooJga6cV+0/P/pQ1p4ShqOUI885Z9/iV60uXAS7avR
Iva7RwRkMkQ86J8p7K/tmlwJTt8t/3p3kfbtN6zMXSZ1FqvSUBkbsbCYTrFSyNU8
jNPOqgXD5Vpbpabc0PtcSEEN/fN9vawGjy3dBOxI2NNR5q707OLiVhFHk1KZnrkR
A94rWyaukD+YIGAILAkDfSgCYuExPUowWAk+LsHj7JK+eARyoCPPs6K7yu0bNRXY
r+G+9WcFN2Lzc2thFJarNsH6roDvrAa9np6Yhdjv2ICCPRTxYSP2ND5FQD9NHl/8
75VwNIfl/kn5p87c1XjIJTPIoIvmIRtICS4qC0mAYseNAgUrgvo3dgkEm5Whmv6x
HqW+E57IKau/WYkBA6ZlILQOUWgC+utdVqxiAZu8CMv4mx2JsFkLv4dCYn93g4eI
nV1tBtBDCPWVXawCa+wGOAH8eLbssevIuhfsXJIU2kRH+rM83GjuuGEeUqmREhF9
thmA3sAxAX4LNxZOO1aShoHcWdD+oqIYE3d9K1FowealoMFf5cTPoIkAQv7C3NEc
QYnmtMyOkoEINqxUOHKee0pkJ20begLx/GJfVtu3MVFs81x6kFluLKbzTd8R3W8d
1eKYAbPPfsfx/upUpBQq/uoQfH8RWwPgU/Ikw8s32r40iiIix5c59VQB7eBbg+EO
cFqxOIWBEFp/yFmuWkAIUE/Xlw0HIy5eSrCAAquzEAxnWxiVUlA+CciXCWYnhDmL
sUn6jFROmfmm504rRDl0SIoJBwJlL92rjEuES+DIy0488/CJU6nhP3l9fhyWT9YG
OKXwnHL5vMc7DH5WCl63ssopakqshfP9IvggDRqph4VuNK8eSOFQ/LiE2o5RHa/Y
JTsip0s+yj8a3rM+M+Mr57WOCWMbVj4Bg9H0VQ/2BgAgO+QLnAAEj1i3J9GkEx0p
j1w2vx0HG3aGSlvX6/f5x1pq9eVDLMAuFMk/ICT/WSF7+PXXIz/Vk9hP1tRgS4YU
IL+Yzw+K3Mn4Ucr1arSSF1sJZgCmoq12/m8+9KnXD2rD4/svjYSLb7IHrqL/i7mG
wvuck+qfTIMknuE3PkjNRtoyOYS5O7pqtbJvT28Xy4f1YTTzaUK4PtbjlQcrMWFG
6EqUChiKeUpK3afbCLQ5jFHEcQLJkzt978p/8uBg87LFTiG+Fy8m/GPqZmrBGI1i
Az3DhlUvueeZhSB3vxJ9BWBztYJXYg2CfcbCrpQiIcCBnk1e2A9lqP6nOW7Lry2u
C9EPHQXz4KpwoW99Vu5B+nkR0GBerO15cWvdZr0UNLPQ0jgcwYTzzT17mHwHWmp5
1tkFVgNsZEuNbV5/wr2FvJSpsBOZpXDRTvRnm0PvTJUqRpNlKRDOul+dmVyVGyu9
Ck/d3imgf+oB9KCa5zsJ9TYR2mNngOAIGu5whLPbjai1gsqnbK9HmQR9buapEyqD
EmUXQQlrdxWZ6Jqyh1/dH7GVOZZtMkbZznNjIEltAMhoes5msJtzRSot9t0uTAfK
3ixj6E8bj6y8Fz/j7zGwS+L8QUX6uM5cx/oli0pyQhvZPzx0NwbD9CgUS7XKNlBk
ra4ps/vbUYdnhVNKoZCZ+p9BRNHHofCd6ZOmaBIvUIa3R96VPw6ts1rarMCqA60s
0Wmilyn2VEY+ut7N1ti7FuSIycS5nwwhZwZbGIFgL4r+Mk8nL73c3NvhC28qmMAH
ftuHbSs6ic3/OM5FoxCgIvxKCogYLS99P8LaTtUsaGwt2IvvrwqHlprZVsvzT/Uk
33B3F82vmKBubBBERmYZqMmCMshhb9FU2Apexkg/d60Zd2CbF+rYjD/dKlVdDRGA
jGqtMEU4I/Tcp00dXjadTVifvdYOb2kY4txlAXUU9FZm3hGJDCbjJirqO9JMJWTB
t3NKjfD7fVkgVWcWzWEi/zdiDMXfBLWzmr+zeZgBUfy5MUeWiGkMVZ7F4hTdEsTw
SdtlkgNS6p1vFxRmX4v3yv9iaCEiEzBg39qF8FKXPWrFh02ugl3jIyAodhmauvr5
+r7pvMB6jOsutpDhpWQIPTa3R4xrfNAWKIORadMgZzSlsDaq06ofnFGK6TNDoNjg
f29q15ipcWS0yc+etdAHXAYdYFDqpW+Cf1UTzY74MmPQm56kXfygsYYbBlBfcFOa
ARQjJMu9dNnAINxA/CaQ4xoBg0LGw/9WrdfB6vjPOzDwERR6YNqFfYQ7cOSIL2Vn
ceJytDsAQjyeHDGn9uBuqqbnynwTdJnKAUz9+HmYiu6S41ag5LWAapkZrTWnfj54
X1rRAHl/Mr+B8xe4qYAoIdhX53k4rzFr63/MXX6fg6rob3cEVptAbas9ut/o7nYS
vahiityOjEcLkuZ3Sua0N1zvGja6y3FHDON5nGCtr1nT8itKf2M5PymtJjf2WxRi
pxK8Mh9DqxbkxJVZCx+DdMbGbCqUVWlS5lSKcZ9ItJWHfFNe6zv4CrB3Tu0gFWdU
10r+gXottcg2MR0aw21VlnHEUwvE2KqIlS6JRKlDqMKD/tmgfAK/5vGqqLYG4Uo6
RUanaymDC+Be+f6TtaqnVy175qYvpc+KALF6b/8SyxdfXPSkS/Y/TqVCvUPhboEI
Qt5U0cM68T9giclDSRfB9WP2iwZIf6cCBKLyVpCuox+SXOU7ZcOEPzo9M3C072vY
nz5v3eNwcAi2r18ZzTbxpe0ctZkpcvzO2W3wnml1yQD+4DqBiX0AbBxHB9L8cbbQ
JueaYYCEZ47XVS05tEl+Po3w20JKWzPM2mFx3zoAC6LwpokU9anVh4cz3AC4/xcv
vbcaqbstw59UbiByOtmakTZJB8n2fm2sGenMMLHer2xqhAhqjjmWuvIjiTYWYrFF
XJ/iuyAS8yqC9ZGG0IvJ01gKQYvzKV0MfQ4aef8Vmz+C8+RVF8O1lsrhiSqjebCk
PhOPEvZOne/nKMGlaPVztSXMOPTIgPDQaWqXN2me+J1Mm1Hj2xL84GovvBj4E7IR
nxo3qwR+5mz0g3MzR9bia8R6ivxCcUUgkGuSgtndNhqjWSivxs9CKuwTc0T3DXW3
U5sTsmrm9NlUQas/hkLgGKBqM2hijrlsW0DoMfx8bcovVt9rFfkbLED4NM5/WLnN
QJElfHJDLZ9LX9Bc/OVe3HvTeijM8GKu+xnw4YjiWeIXr5EztvWScztAef1wLn7W
ifZ7MkiFI7vIkNKzw7WFow9MBchM/RvxhYfl1Mgycux5N941vNC7P8PWFnP+xohY
/CFmyhPiHEufVz43wfMwbvfVfxLhLgkcKdtYr9VJ5EeuF0oBcXXMwNlDniIr3HsY
tijLPJ64dC/jtfeNOVx0kHUh5FDaN8k9PKAyjuM9ObOLDAcbb5RswTbCEfrloaNe
HCyrAKUB9Omi9FXkIThTlMptKDwO2BwGbHqFMGfw1kmvaHYVzu0gcM5tACy04RGL
vXwbaR2LfPNNL55Dq7b6wat+d09Yk9bMpQZcIbgvq8oBDEHSL/wHQkjuVPPjB80w
E93ng/Lgj5mEBo8OMyDoBvUMGQQNnrnn9jAeldueusqowCKyglrKZoO5V0kS+1kN
nSEap3YkIj+/1Qy5/8e2Zvmf7D1I7vi9SziQCPMEXZhXGzlzXT7QNkHz3xsyGLx9
V8gOHGzFLOlkpHWmTLci2/VUhYJ15qmLKqQwk05V8Wbh+uyRsj4Mr86liQFsrDDp
tUNFjPoQnBE8ujHjloXRdQQIfIFC9DYdCto15ZQ7lo/zwgWfTW1wviaxNRmtya1B
mtwQBJmJDlmqy7bY5Oy8NJo2xsFnBduF7wzuo1ALvWxb2nTx96H5sNOgVTA+jXQn
RC9Oj5Jxx4t3aYXQO8e6KHn7Y3HJ7OutOx10Eqa6VnnHUY0rfn+MEnFJ0aN9P7t5
9VLkGgkBlCmQoxse5QzCNa1VroaEyXSORzdbZnpjS1B4XiCyy59Z3clvmaWU9MOi
D+NjezErKdTuTnX0zU1lKgB+0uHc0ZwIdhSNZFB4uzLtTxOk4A1tpCMkVX2jzxGm
D6120qLxofmPoOaQRtCvDlx0Nk50BlaqxBoL6QddRGrh/cR2ZjXILSwl9v8Cabxy
/+OhvOe9hIbpVt8O0iJRFxY/vKrmO54uZ1jGOjuFpLTIsYKnMtgCMPkxOZuBmwGf
Nqv1hkCwawB3Oga+G+4rwQ+BQHTm1WrfIETRNXchFFB5anbIOjxS095BAH33Mb4L
JHwO63lLotlWJs2FADXVrUrpnFrH73Uk6vznMEDwSDV+T54WIWA0AtC1SCSxPmGq
jR3xxK8OoUQ6oHT4H2L23tl2mKBU3KgCla+yue4lbmqr81oRPlJM7ZfBMqG8xtaJ
6JeAw4nVAAcrJTgtfFiaegNXCZKs4g7ZVL71MNAGQxAUL5Wcpqj0xtEj8Zx+PoQm
B3k4UsRL14PiJcNH52lZ43yNdnCpw9j3qxXH/rUxF9aOJE1KZE4EfSnaBZAd8wzf
JhvLEeXZmq76QVirpKw3fPwusSOJhwNVIRXUqIPJV539Nn4VtDxb1kaEaxIVuQEE
oYtS3cwJdPwuH5QJ8uLlgyyLxzSF1SGeqpdhvCvIZnwIMr4sEn8YsNlaKgk/eVQd
/0z13iw5CBm4fdg7EtkjMVxGv8MEmuoqPh+2NK2F2bciBXXDrhT3hOMqnGUVNRhz
KPzDcRViNBqiFJbb2YrH1CcpkKbn9og5HUFIg+fXexFG9DpXdwtqrGZg+cGiqS+G
f8+b1RxDtxIv2s2FvAhk/ZOSFr81yPEBERQX/yH02SUrPs9XaC5W7PliZ1xivMS7
KfK0egENdM1Nj3rxgrPQDmAt9J73yTycag/8e8wc9HRCsxASdowZ3sBZt//I9/u/
n5kJ164xWZAJVxQdr+kqa9tpHxS9HxlBTpbCU+RTRtcoy6jBhrIe+DJr/aZKizik
+E4au9frHRterRTPTngZ8m9nvQxDKJX9LZvyeXhRGHwFEb7ykWK+hRT7XHkUgeR1
6Eop4oznGyoc2gjh6dXl2/zRHQpQ/amjwf4Y4wNDDjJga5T/oPc4oEaVcr2xRypI
tdYYu5SF/qbhiFWy8kE3qaFGIXOKRDNqHh/qA7KYTwlsWOaQ7WDLNnxBA9u3Dgz3
83sVqWmvDkYHh1+4NqoFfjE5lOdVPFHo4rpY3QajCbA4Suz3tTqF1Jjye4dBzxOL
tC3HEPt4zzPjbxgBrN53O/gcvpHvGE0GO7lUNnnL2cgnIR2acnv+YX7TQIuEHrFs
NvsVtTJSp9/BFSH4SdgDafs6oAibbvmZoim6rFJsnv1X2driNLSGT/4T22ptC2x/
0yEytLIj3CIq6fczqtlIjqxVRGfU/YAhhTMTEntI6qEJjCpWbBPlMVXH/V9E2Q5t
RIj73FaE6+Mkaf7gN7Wdz1ZJjTL/0RuLIUn9+EHkKUpHOFHiHN3VSvrN9dpWzQNK
8u47IqXQxYibyNDxpE4ksHH467Ft6qA/NagDX3SoRkTglp8sc5Ay7tZJLk17ptjF
/Y/lqfrWl5PayXwPqtoRoD3lehn3NKqyhdDm5v1vik7PMjkwNBrXY6dbYfk93H22
Q3h3La5VXwr/rddfvmIbhTrlTUwnJORRFD3SMB4ZlEePEzdrkSv5KSdZf9UF3v5u
WsWBsdDT14LZs0MNOrA8ywIczTOA+Eq63F+coq8y3rGTUlhvuSsQGlZ66zyv9Sfy
1hTdLVVlKdwgQwOFJFHygSOKfUPwMfLOicRQtD1ZyNIPJSWnr2muNdnnlDkm34R/
1NYcIqVjyI3DO1fW8im/vXNNsZj4k5mdQ6STATCB1LWP8P2oYIZmOeXcL3YrvD0O
/Fb/ma3ZwdHtu0ZW8siQ9wd/kiKCcZPXkjA5s4Ah4c0frhiwSXvPPHXEYg020bTJ
pc8x2O/KbWE72Zi7lZm6fRkQjoDFRIKw9Mxfy+DCoxaixQ7uXXEwU6XUhLGnjmsM
YawbbFEBkXd3p94IVSmq9zB3bFRTA6hq7ZKuCvLL0UJHM9U2gTfPGW5Zo8GiGJ98
sjAwkRae13Hj+kN/16c1XzetS/OuS+Cb8yhTXTuAhJEhCgZKwVlbO3Zvq03N3yPL
xGsJtkXz8+E4ptMcwPFC6NRJeyWHd9z9GvvOyFZU18FYcLTBzDstVrc+s3lcpQFN
zZmmBCacTJC15LI0VvGpECB35GqPmGnSd2sGXj7src6Jv1IS24ufDcxIjGq3Ff1o
37tNJQpWY6HSO4+Xnt4jTiv6Y/7n8BvrUj+VMyIAuFMkKp+RfNCv++3/yY9Jvn9r
OS8dEU070yLaI+tCiFxpS3D37aGibHEDM4K4L/2WgUaQKWIymLnIt/QtMfFtARvJ
Af7LGMpKzZC/zc7NZZ3V2M5fdqPpvBEqAOJUFYCqr++I0HyiLK6mNc/g0u8G+v3w
+mMudZO0KTtFNwfBV0LoVIku+y/hxnOcS/JF0jqEzrSuAcnlMn0If0TyFCpffmBH
UTMlP7VVyKE1v/GC3h9oiA6o4AfuB3myTfPLHupVjZk26YR3dPcyIq5semW9cBEj
FHtD5mF2VypxkmA6n9xeZwGc5KW0y8O0/DZbGaNCz+LQoetMrD3fA0gBo5wJBVMH
DQN231rCGmIwT2PYTb9F6FhKzEzD2ZlWLJkf1P3JZJKI2W7TBR2CeL14hFIApcY5
JIq1pdFhRuxNzYxuIxLuACBTwSaFWQGGMgK6SrLfr+4UjMj12c8DqHC+WzEJVrzy
Ln4A4m7QWSwi2Y8cNgBHCMY1OSg5VQ3UXOzcB5cLH/3ybuFxfbuM0LP01moSRB0X
YTjg+MLVTIMLZTfY3TmUiTol3YBkZAQoU6C0ANqNxQ9xc/eHv6X/0PQON43PYO7h
/OUC4Xq0tiQXkBk2+3G8FWYE29pbTpnk4rT9N/13wunUjRSMLh8fE5B9LKmUPlmQ
gnaEAq0jAxeORUdC/u6odTJe3VkSFJq25ag6c10tbCi/03M0r+y0Ytf8h6ueqBwj
3JGcrAkrp6XYc7imbGrIZy129ot+FPsNn9ReapgCJyi72XvtoDvd9Gfv/Aidop/g
gNp8mSvNQZE8aKsu4eMiEfF4NW+0IBHtSpbIzNssZ/LDUvzSUS5O2nvQ9MJMdcqB
tUrifHqyh85FRB1fMeD66aBrn3sp0ioUzAhmdhHtkBiSHpNA5MaL9edHlq+GXbL1
rC7nYRhcDbPWUy8GpNsrHP2XPCzy8FfvUzhmg5TkPSrkcSBb/JK3uN4a6d7HYoVj
89NEeCrXo6n0twPBhvx/dMVqChuH4mRhlx+sgSk3651s1UIeCIDhko45OiVF4K1r
X6FTsAgMZtIMyM0iYmy8jgnIOx56IrOmZBZiGekv6ouhkV/+PouK8vkXFltyViQY
ol7bFLiF6fsxYSkNjhzI4z39L3yISbt0+lwREmETNyg22xi8eRdGuzUYP206izAr
xFoJyYQMx6PuFTSTHTx4qRcWJKtuDNb4atKzlsm/E2OjCex6FEg+LTD1ReCciiOQ
iqtka9MRUQ7wrUdSAD37rmw8rJW1MCUxYzCQJ8R8YMrrLmWD/+xFUVXpbA+dOxhE
YSY62/BmuyT/7MH+9cO+VYIBD3r647ZwnatcBudFinXrbC0H2blq/F4h4P53qEKn
0JS2dF1oIco3li7k7UH45aWKkQrcXafYyTRgRFIFoVm6MSuGPe60ycNQx9U7FMG8
p8xvOwjT6M3KGVChzn3u2zLuJDLr1/Y6uic3xwwMe+kSEHtBzRuf3C2sBIejm4TC
HLdnIf+CpA/pSJT2j52/7KneAdBt7rBrDZzEviJF0TfOcJeC5NkFBzFsdVRZuG1K
RoFJ3nBe+YTj4q8Y+mXg9KwJQUoyp7LLhVLKJmddcNaTQsd2WK6MM/7VjlkMK1UH
3nxvv+toB0CxuhJCWQIJxIoJVNJkX6bY/lREB6qfNwUqy8R7ip/0Yz+DXMx+F9ut
a+oynYoLmsM+yQHYN5OJpPIRbeY1qIYzguvtML7HnIVEFcODQ91hzEhWhTtw3coP
NSUJfkahPmi9x7yP1cHxLZQOkEiRfTGoIa7e8c3qm63Q4YK3bfWLntSv4gcuDnUY
xteok+I6NEyoSoTDAekv26ooHcJklEoaS2AglihYQ6n0252AYi3+ol5lDLCuSdje
EY/mV9UphRihyTlCXQ8gY+M/+ArNoxhB7Bo3+2e4O+mjMqLrQnr0M4Dn+xgVl7cQ
kTimrL0GLIU1maZ9JipK0h89bEBQqZWQ5GF/YVQnLLfvFvPZ9IR/GZK6/X9goeKf
QUCzOZGT/W+ErMUfn/cRHg+h3CqOcdvqfsq12fMexO3aNSxH0AZuHOHW0bWp66EB
TsZBwB5kiAQlA04DwfJmKUWNN9JbmY7NREyKjKcAxl6B+QaDG2GDkSHGfmdmtXdy
M1BrSVGYT8Ka/H2pUbyyJEvx/Udfww59l2v4posxvyDso/RzSaXV3Z8JmdlZDFK5
lHWcr0Xpb883pqdR7e9Q4Vvcc7UCAWzi531g67eScGhmFqmAcmY/+kWGL/hytorq
o0DysMWpTRPzEqC9/oeDtI8DsN41yDH2+6R0DAK+Vl9Q50AqzpL8NqjPQxr/bp+m
3Geka18afTr21lTV/nflREzuzIhtgjdW8Wrc1jZDzEag0QoaF7ms6OmZSSY2qS4+
hR6Y4Jkt/YP88htu7YrOhIv79Bli0MJJSLkdUhNsQATAARO10IyJRs7nhGSCZbIy
TbQ2cUhtCpcUONOlxSM81zIPptr7jmS239kDrEymz3qhZfYHDAHwTkDo9dS074ij
HbZpheYKu/O3FHYFP1fVHfvcKSo8z3FG5noO4KKaeiSPQEsZpHWRqFQ/CmG1K6Zf
8waBmaocolywDr0cOD73QjwYGwnNO4V9q5XAe2LVBYdPAt60Spmm/MWZuJaOgLmk
5t80XsMAHtvQRRp/bRCq4MYhun6Ped76Sb845zq4N5hJw7boQa1GoUCuy0lU25bG
pxGxvXN60I5GNM/4sf/4ypBBuMSN8eH+OgbvznUz7acYrKXBwvicF++UkoLK29BQ
S3LO7K3J1SmHFgTbGHIjWI3k+b15czUcUq0qDloDKQmCQcKkAC0gXYpV7p3fmgU4
u9TjC1Y4N21QHfSCyYbVM3BGL7xfq6wkkVNQiQarrPAUWlVNxOeqzJFrxPhRZUxE
RMAp4RTRQUVqEgNcsTmNfnTt5ehC5ErxnrQf6KifHYcaVK7OYZebgaiFuLlpKes3
SdEspwMFCBS5bGAi6DLKrEPGwlMh9/FC2paK7P5hd5hqHgMNya8FkAEtgxo0i3us
oEmamudrv5ApTDnFBACF022gqcV2x27G2QleaijvA3MAsA6R8dfAFXsv2F1XP1KH
HFsqKj/zI4jZRoF95sJ9tIVrlBzWPMQyIC2opWA7NZsuCT0f6Hz4PvUaLJj145f/
znrFoo2b6vU62h5FLLMY3+blKFovtMeFuAKGmogghvG2NvqsX7OnEEMaYMCIT6HA
WgG4OgUnhMXZngnnxo2VycLU3cxPUGQVqvIC+t/+Zx96pTBCSUqAduXSAIdvQDT4
Scoo+0UBK+k7s+Q9G65dGzTqwb47JpiOIAhxISdX+aF6xVZXaOMydkmRYv6aKBXC
D2xyVg4pqFDJV3wKe18C7oTpMwIS2vZse+D2uBjjNpHfqMXHPQfXl44vfT6XzjZN
vhG7/Ec83+eyfSnjZVT8RvALhoz2XuMRbUfWYqT/OG6si/35Xuyj+Rngsz6ZVYyb
PW6lhks/t2iTEankJR9iHP92ph8jWBsX+uYHhyurthguVPniWl1Vt6SuTIB/IcpW
CJTZ/ia9gXXOKSLDR3YQTMXlK7z6tF+nFAgv6QML5qKPpWSESRloiYXvduDQOiy5
HwixGobNjD7ePkVokIMg5vSya5qtxpRGNhPAAsf+vdjLzPg4giQeuy+SI1bO5fDf
7oKK/flalsV69P3WJRo/jaSVql6JtnKNnp0kn5miP5drGyR71tYOSIiyuAGXCjct
kzGP3c/f1LMaRJoJ/eDpste5qILUyhgTsdqDtyuDWwqiGg5iOQ1NwT/M+1Aaosjg
DFjwAeMYWXbAQXawdnaF8JlQLYl++emQ77Wh/Kax/CABybTn+qyIJJu0/mJdmKrD
hvUdvzjkGjmITMmgvwH1nXr9V6sAGt6F5kYl2bo7ZDt2ms5RTuiEFBs511i9rBAM
Fu1+OyIH6KkBkddf4xHZizK4t7ZzyGTKBXIebgozneLPc0vZcm8RW83erHDdcBtQ
Xrj3/o7ynnATGfgEK60NQugYGq49Xl+wcKOsKGq6jN83BxL8DEXt1IsbomjTt1aH
didQvotpwfzW6JmE3dDgLWpKm+HuBsJ51KpBNzpuguoAdqu8iwQfLrLYTx2bB/wa
spGUtO45sGF+qn/NM8S61JenyOaWuyP0NlP7CfRlKCR+fnL2j99mNswL2a8iBwUi
iekufTdeyl0P9tOsqs2SMhvKj7p964eNrJmF28ECrzvJJsYNJZPm4MDBMEvLr18d
JUOsDa4qyf23Qvok8uNAln+9k3XtQUOzgs46OqoV6Glc7UOsWh5YOnp7xYaK6Lau
wBrKBWCbd/MlJgvrY/kUvPqTyqgha8nN3Mp/PnTrBBJu5dUFZtiLa0W+Ib1gmrrr
S1n0HoGAopiULy0cCyJG55S7z+cvFuC4VQTCxspeMmM+VCG/+9KEKbYMBaTjFFow
OgGiBzABTFa3BAOn7dtpBPZVATvzzIE92PFBUZrPKPUms4nOET4d/dVwhhkGAzpq
mKNDMsFt6KhXIUF3Z6IkFRo7GK0OmCO7wG8xa2e7BbZ/UyWqTNrgR5+inaNsL9zO
nGhnvti/J41UEEkXtIG0QqqmivHy3vBx7GZJ4dV39/SdNNnDQ8wUTK7SOnu5/Xr3
zwXADkul5kCKloeXyAGP7rWg62fUjNx+eCgVk2dPoyyXDDTgR9K6cJCD9PUcQkda
c53qtl8xKNhQXXxQ2ig4IqpAIMU4Qe23KfQtGJ7frpKHQM3h6pn5S5NQRXRNiIUZ
tJEg4hYZETeOhBFNb9z2+N/XwHve9xj72Ob7uTFT7UznDob3JPawkM6jOgp6zH3i
xvjnSBejM4FoCr160a2UZiqf8EkSYfAlxx3CvZE4fuCZu6htChAi0usobBYQMUBp
2iTVnTL+2thgjEMI6Qjiu7AG78z5+hU42t0qe+esXMA5LJyv5ILL0lFhbQqTFE9D
qIj5o1MepV+6QO5I5ahML1cMSKl9G8qBttXyFWP/CfdTT/QACGv+Z7GJl2scUGof
GpZ4j2wyOQ7tn0CAZ5EuhQFXiLoMXa/07/7tAvl7IIR6tpbyUtwFKbrA5JaxgVaG
yKB56UqqwsmRkC0IjWZiziEHyrt6bgdks4CkKaYObwoud40N+wlR5iJL6WmT2Mh5
9mTtPBexyEQXoTsSe8MkvU3NpmGIPmPze/DIDABBgzgrRdrhoBjT25/NwSLmhZNq
B+H2BLcpJVXnaSL5ysjE9LwDvP0ksa9sARhBg8KVkwU6JCltNDcp/pIRYy9W/y6w
25SJxSvn/gDevT35L60TNYvOi/uL3bzG/WC7930iVOB+7lK6+Hf5JGfafntTfEOI
hNRUJUe7dQiAxajZrcDYSguOJ/F44nxJIQhoOl7cmHp+d5b8QME1A/OTwZ87cgi9
NvrXznW86fqOejinzzm1hLXm41w2UIHBT3dEHvv8c7W1m2sGAUlKuOE5tQGsvqw8
FLPUVatIfND6RkM5blIJyWWAZs96snKut4lhQAonD21xn+xwjuUniW4h5X2o5eLI
hAzl3nhKgs88glG2rGmCHKVtV0NBQoySVi94f7WCbtKtywpNiJDf/byA2EdR3BZ8
p7uFV/kL4dvg3CGdBm+0LENnWDvfrTbKlQREodpws3cHqouOHbI2EbCm8JmswwUX
K2DJ7CtUw3fRI/3kK2LaCnb8jD/WdunWRL2efFrvMat0Eoz+wscOW15IAmKBcKT4
PW9kdhKV1ZITBEmRhOcGahcJvf8arliiQyb9ArhlsxCP88gl0SPg2LvzkcIelaGG
m2TOhplUBRelg7U64l6yswBwfK8Sn7C1K5FLqzXRxlRMISDqozN9DRhfO/iBP81e
mdfZojuzeNzL+a5upSKuvvYHzraqzn2SYToT4l7RkRDXjWhEtJuuwjlS5AXYpx7U
6smm5AfVauEytlGAR9wSn1RsChCsKLQHoDk4IluJNNz8yfkN+Ll2/ue6NwApcojF
oAr/rpZPX+qRp+RDk5i98XCP9MB4W9ZuY9+jUYaiZgT/h8iC7gZmmsc1EZbdvN49
5m4GOeycEKIHx6OxLC7CBU+cSJnPngLCNRcGyDuhzbUAjN/8S9Wxf7Z4ux5ZT85h
uUSJ/K0uBfqcQ6caLZ54jhyGEnARxPdURJ8kROptrH9j8BZarKDKWNidwmt7aAG0
ftusqyCkUQQsRoc6j0BS8WvV4ze/DJFBHlnzpqxUGhtOjro+QV2D2FMopN+ExIOy
vK39BioVQOqSHxr5RLkR+pDgFSzZ0DRjeJPmcWDpLipnTckQwUbfRZdd0FnRffeB
dF/3vCMDEwSbMctjnMT5XQMqNuK4f3zQQ7456zxZjZTKobr1cg/7tPGE7N5NBPIA
8+76o0x9wohmfn0LEaRYjTOqy9BlsA6nFr8lVPcFl2DSLdsQl6Y1NyJPK4fFdHZi
svIU/78Oa9z4e35PzAn+Lpl4pCtTUAL24La6L0XDADDAW23q7XO5fh/CPphgHQpj
2/FycqbLvpZ1Pe7Gh5wLEI8UhzoDZdFYBtPub0KktZvFMPtr8kOrtgIWOl+t9W3M
o0Se2w63krHvGK8CgYxEjbQhlBf9dTYdLdjeLuf2FAPZwwx8uzmN7JQZcU5rYcAk
IfzRBeNGXfEnp8dz6aNVbrXADdjKe9w11znsUdzJRJPB3bS/Z256DyVatFD0/eQK
zFidhcaoyIYRqwAe2AZQF63MX1bIXNzQDd8oE+C/Hu57Wv9ennq1NO2xCNjB1hAA
lWzasLwtS+Z8t2yuoF5Bz75WKRJzH2KEoV2j7NLdON4RYCqVIqQ1JxCpYEcFyqPs
clBaAbXMhqDyKaNaGj2CSev7lALjnV/HOl9XQB0F9bog2Y8jy3IS1y1rgHFhQk79
9yOkRsKc83ZqBjh0PqJJfjV5x4abJNJsZd6p2mGFBMZEz3U4puJZr4lzlIKU91mZ
DG1okhVZWr7+QS/BHxQTMRqSQCXRGqemgBtsiebTUToP+e8xwk9j4JHLq0CCeqaQ
xVpZQqTf7A6G7PLNGBWMsh5YetdI/WqxMIp4Vjc/S6bqJW4sTVzwPYVdwdETYNIm
zvYjNxggRYvP+UtMikQWg06P76Bv1yGR4vC9STIFiPFU7vm0aCccd309EqaNqUb1
zFRBMRxJPYAysvS2CFv0WLoE63gRnwLMAmx0NBH9wJapkkvSipp7TABTQkPXy7RY
T5UZ6p3L8XLjbTkXgCKSfzctGastDaRcjomqiik/qrx49xOF3sGYALAxetv+jDbG
1dlvjmnOoE6ZcEmtyjSX2QvfOkRV/cikbdzhom62oVmrESqOQwHUNUvtXk4mNlWQ
0FfDL115/y1d+LIZgJBUUXSk/i0FFUJeRipaWMlqRylUrIO1w46zu5ZmVuThufzU
tMMZbrNZCHrOLmCfOTq8byiZBbTxT83+gTVNPq7qzxJ9rqyFeGiWIxSqhuPLNu62
KgeC9R184/9GUDaDjFsjvWVSib6wCzRhZnY5CPbZbq5l2gxWafFWWH+Zv7v6FdAd
/FzfxpuH4n4tvxguQv87N+UDKOEMnkUFfd6dVamGs7er+7y0akAcRdsoSUNP3wxT
aSHdbWrsrAcBlASbRqqd3SYoUDICLKMfl9THq2OMOdtZpc2CwPOLNKcQg504f6hg
YyS5m3ouYsORQgXFXJqLYeONK9o2GrMi8kiR3z7fFI56uU2wRpYmx3cfQ+K3M70D
ExGy+NQ6FK+hsrBypw5TyS/gNw53qxFMtbQuU4bSrY4/uU+tD9d3AALANh1M7VOq
cIC73J4eGr23co1naAJyTzS/mxOV2GerPJhEa4TjwkI3znIRlBKi1O80N6i+Dzqq
0gRg9hHuSCn57hAP+jK2UoQcZ999SQuiBk+8v8CKd9g2aQz5UuH7TdcgLEjUdtJN
5bVdt70o2YBtehuPPM+AfMe6TlfsOqEUpiYcr/WtMcsjpn9FfkcAxSOIQX+13j5q
dTswrnrqeX97iSAceaGzJ/xYjDvM2IgDBZaDEzcCdneQv6o2mL/hIfyIZqn1xLOt
ZCG0QcLM4pgs2xUsJehwd+YBeCWWfSwkIC6UknIgU5cO8g1FRkfOqTP+y3Rkj/qw
sQxc31iqM+8aNjCJkPnpnmKcknIvEoutnZME2uS3vMgnJvvpHqbj3fAblEZMMHNk
fZ2PWSZU1jbVn9UdkfGSeywk498nI7Rp/Gq5cqDpWXa5m/NPonbKnyclUJ0xQ5fv
W8iZyzKtyo5M4eEsPcpFWVSPfXPwjrCzxY8oYJekk5V2kMyPSweiF2fQ/6EZqcmB
7ivRvHniriLeL+7CNlNYIlLJudVx8cSYnNbirpcCHvPSTfxvlJqq0LCELSgUjv8X
s6RY2AAWWcN1O2nSyWIoZpfwcXAhK/MMKOzYXouH0DtLYot8m9U6Re4TOFftObCZ
eIuCS2qIq3n0TXbZ3cGDYAiyBnIgBqBrOJubWXz7aVAs30d/mV5W6bX1SDKACpa0
+wJPETs0Br1ZoMA7ft5U0ueWO/IQ/ZmbZxau5sXMEc9rjy0rFO8Fy0icC7Eq9DnR
/xE/cN9aT9hVpI9pdgkthDbddzmRmziidcByro8o6ecuMfr7Nc2UzrDBwN9mDrUw
AkYRGNGdKhmJkueFZuvyYyOBp611NB9M33IR57lTKVa9wuRFdhoIOgNpz5xx3qjE
jwcczJh5o/jPM5CX09iRVdTFDZMbSjNb8m7JTFb8zJd6Gj8+LsnibsWIM0b+xPAq
Ofi6LrlHVU2SsxWd/n2rMtm7SuiboLUCGJH2mwVtVhqlk1TQj1Tp7Qk/aOxSH06u
o1Ff4BT+hRcQpCkfz5ZjxS2VjzLr28CZyq1HLCIfpotk4AUB0yjAdGYNBNTdyIPQ
b2CVoSQ4dO2RvI615xW/05iKuQIjODJom65xQz5AV59SACSXIKg4jUgGZ+XAvLWl
yolmHJyldasjm+TxahbOPrNd4RRl+mJiEBXq80ixh4c0WXl/TIrFM/8ImupxbBBI
0MPeYZaUqVxbY7wWl9FxivFXzLvYQjnVdVGgcowojjO+ZLf5aaFA/Z4nM/DWIvsC
v8cht7VKAsG2Ftkz932igbRCI/2Lww8romRQLD5Qoc4YkSGckTPMJb5YPXFoHLft
ZNW9s8yVgYxo3zfgS436ylTrgXGJqd4y1ScG8xKPyxwV0gOBwNIixNJF2BGHHHcI
KgzSc6Tbl4rD/5i/cnsnl5dFhc4sNldoQF7VXLmgYTqoBT1hn8QmBRtMv88yP1Gb
N0fJU+rBU4znSew73U+dOndpXbBaXrkkIgprD5bmNswBjP0LBglrSrDhGx8K0yp7
Gonu3x7ulNN9uUvn9y5aZ6iL/CC+xZduOi4Q6OtfifVvTerZDX3YJjdBEMTbNMRi
461/7LiwYo6jm26XG/qy05OwrIpomyv79UuM7nL9tA2H+3PsO6cI7gKO2bD/60AV
hGijwkGOlOhpLEV+N4MyQTFXNZkLE79ucTFJjGNVhXsTx1RayvfHE2vPFZeOxQje
EqXoRGK0xFMo6uCyAA6rWFJMTkvAxni5ZP3c9rjgbtPILVMdrHWpKVpr55Utkq6O
abT4GQWbL/7YytMye2JkXKExW0bag9Is8FScmWXTzK+KznkWAe9vvwwMayscGviA
rw851SXzQQbdVLIiwGRRQKxY2+2VzPpYBFrPs3td0FmSshyamOeW0UBULgtK17c4
trHYbb3lXyrghiylTflqNQhlcUMHnI6tzDsSozG52OU4UxEmfQ4d/ftFdvjZF3eE
Pu0jfpf/O3o/qfSkmky/zOpZ+hPn92tEcOtcuXhUUjal3AFd9UXCkDY0Jcp3rhnt
tvcH72+H/v7IZLfSOwLTAcAW9ygdEJ3JG8OxdF1P45hpusb/CXfyT0G0vLwBXGeg
wwQHHWfkid+5LQ4rRW7veV86CRyZ0m/fZ4WwMeAinPA72/aJZuQc4p+zog/bJUbN
djMCsQZqGO7NhQNrlGlAtNfU/+nZPtwij0u59RkVpwdhT8pNVxmvBIUjcQgJb2E1
pPMWM8/m/OHXlyGpw0apwDtwp1q34Phmqg1EUIFNLX/j8MXk+gfGwEH5sVlCI5Vr
UOIb2kG+2WXFDpN9TldgTuh2qfzSPI4nfCfD0VfJcs10fLndYzPGU5NvwhHrnRDw
1mCQUnEjylgPmwiU8hpkcN9q5D1nn3xRA7/d14P4vENgItyk3h/gA2YAQcbXtMJ6
iFhXhrVg8jUTkBN5DZ2vxgj43ICJhgrH3YKCU8T2ZWjy0QUJYqv3Wsk45aQt6LOu
nnfNll5IfmB3wp34oQlnC7Gd0QrEhUhj/vfv2NBKLaGONkPXEEozVxzs8fwMIBoi
LQtfIBAj9oD/eSvQyGtwCa0PAy+3Bll+S8My+4jw8H0CHZejEopyVjkeUER12uNj
st2HK5qyWlKbjR6oYDGczESBELjQFA4SxyojntXL//8vcLXkuPILqteCt1jr4Sm0
Yr11Ac13o06x/ZV8REWogNdC2eBFxG9O4Z/QoziegrZh7jyNtDLrBhAyaNjVQv3z
lU0N/HphCJxEAstgikGZhLL2WLWDlD83P9PRJZpWhW57g1hhTCzn26ajxP/wyWBH
HdApOvI3P48B3+btSikCUww9QbyMgpXvWubLJVsm2kcrWCy8RDj20dNn9AWZnpWV
e8ahnqN3PNCiQhJOz1zzocDrNtuJ4I8GCkeKQpBCrdCSFZTdtadecnOJEUJXBtka
uzt30d52shFMVIszmTaYwpDoN8n3p4WKiXYHqgCCKouep/ibbAjuxYMQSLP4gNMl
E2mm7e/p9utgIsUw5+M815vk4f4eMA4UPK5XJP/33qhu0U0MT9B8034pS14AOPGU
NJHfoKZf1zeyDP+81TdRxiOlhsQUb9lD3dMq+1vwCSvd1kya3AEAZUGkv0FB9Hl9
FmfaeBazmdfJOeadwsOwhmqeq7vUdlUj4CNsEfcpjGzOCJjGWAFzQ+IojicEryA4
3JcKtCXIPb1LYJChXrT4AGRGzzYKJGs5zD1Lx61PZYrwWX6zvVEqqALPuIFGmhP6
onhVHVW+MEwR06l5+NNNYLXpQw/f4MCeK2uy8lLxEXJL2qyoq2YmK2uIyIui/kF2
VZ5qHsxloseL+cw1XKDKEZLaFX0WDRy/dy/QE+TBPiPG30KKBd2yVeZjFyFjcm0O
EAoJoaXy86LgKwxkJ3OvcaQsNb5b2c5U47pUW4Z74Oas69oa8wgcuQRK6w5J9i70
9y3y+kRyj1kBOY9sfJNBr7DFx+rD8FGOj4IEeq+YZjuMBWrzpwitaNbpTghzugIR
giEvxaRgTfRgt2D/CH3gTuyby6HyIHsWcGcEtlLCAjRLjcxAga5+C2hr489sw1o+
XWMZtcN0x6jr7j+Jor3Qqq+/UK6SN7oJP5CKRb0HwUiF5PxsafBrIyrEk1KvyJbW
XKnN2VvVjcbUdeBYfZR6EG+vw0oawsPi2nH0FW4s1FkqZI79yhRx5kBnPctYNQPc
GcwMnktd7wq41tjPnihYoQfJ/dicefkuJtZ44A9hXVvI9ZoT7gHbdo8WlShOdm97
7rJowOF+TbXgUDJOunS9p8RIiHthnMCOnbanDFnl/fcRHMTYqM9n5HQOm4leqxa2
Xswr9ZkxbAKFjRVPGRDNU5Ij76dtJ51pbL0QT/Bw+Vee/Gai2Mv5nj+VIxsnyuFP
uU0lODLFt0PrAKgN6mMmYCvfXcdnmO9p0jUxJX3pjLGxYaqh/3qbOU++4fm2ak7H
Z5oCwqqNW75cHqCPnw6tPCS8YCkM8ycjg1VRhAKz3nv3wfdcqb0MXBku4tHDA+LN
yBhLnxoJFB6/Rc0y9RU+yv5s1bLV3WSOAsSeSCr1mvh0O9Jw//RHLa2DrjAQhxvB
yY1VmSbMOxxiJUK2kRf8HnCkZqnGbo+9A54WAHSKs93k4YOgWkCQBVALbD/iEp9t
6/otG9/IqjQN5tc1Si+MKy9BMH6H/Tt0lV0y7RN4GeDsXG4ORtlUv7V6PlfidZd0
+YezoFgnGGFd8u/wqtt9qlFTVsZR2mGkf9zrfbE5ecOeOp6xYuGcpLyhduzaUwUM
BUUjve3d/6Z0MYi9L0WuAA==
`pragma protect end_protected
