// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:16 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kdEPT0fb6sLTxMVW5q1ggQrigNecE4U5v/QG+sHHFmRflkMtz9epeyX8iukFni3S
x5EuWulVRNyQQo+/w6u1QqZwrgmajEZNPwZd+fMTPaYMGpVwcBcrtJ8jPt2fiSzj
h8Yvr+KIJ7lsTszKONNzX9Q1JQz30j0xQ4rNYJ3XrG0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
v0fZkwJNvbX6Q0CCir6jXClFxyb7mGHEIyd9kRx0BxcR33Jf7nQDInsvhtSOZP0q
XjxqCzFNhdMO2+2xvVXPoTxVO0DP8SzHM5KlbbPXiHFVr+FqHZza4ow7kBVOLo1F
S9VNS7K6uq9ngtD9fLKF0xlcaBcNOfRRqQJs2RyenqtrpXhWAl6XXj21LFNFiMtJ
iYhKbTfxgJ9em4Lc6LHAaCIpXt4FCtLAjo82LHJwaAgIm6/jP5Gf2xByH5CxNtih
6bPbwkgy2W1Hvl1Z4Zwpbk/aOqaQ55i1ZxVhyf0AWvg+Olvd47Vweyq/C4KtjZeJ
tm39cN4HNzq/elqirGLAMS1B4FAxp93a0fuKG+nhtIsChUSbqi5zZqDrUqHNGuMY
xDB+3tUJHTgL04JC+5QmrtWsoplcbPqJBHyygkCnrge+DmcPZQrPl1r5+OygUM6I
C1zlk431Gv1t51VWv4doHniPBZgt6k2jSdR1henR5q9wcNr+kwNfClPlCa2wBLyJ
fyGDBe/ywpYO5HTvzlGNsj2qQ906habfSIW/Mq6t0ng/TxWZYH7mFWPwNpJgSKpY
PdcG2MlrcU+LMPDHS1yv83FDWgTR9WuldhMBLsTzXvEQ/ViWrvsHqpM2cKuR6ftB
FunBX1Yaj/nUuR7MRTZp/qAwEWSlGtsgvPL1ZHgekZR/VLGQw1/noynXCj+cE2k7
LPJcjWX5wuhpxW3LjXR1zhnkbr4FKaXPnhfPaQdW5uyzweXWOxjbEh9+ZYtYOU2y
+f4RGMs1ZbDPV3w9tUyV28fDRB3i3fQWB8GYqTbXlvUOGwiGebLvOGuKX9sK+dxe
mdIazTbGfZMSNxfvTSe0Lv9JEnY1wFssMAeBmKg87HPy0E4t/FTdq/UXGItetBuU
9sUhvjjvQQ9UdIFX5u5RvHvWiAE7TTBFViZKKLESB1ibmIzl/+g+MiOUCbWMnN4W
8CFZSFrUHpPJRypkMimkSSjrCZNV5jzrUp1uPvaoMjaF2Hp6yA4GMjjPZldEQ+TY
BkCkNeClIeOJUuW2O2uoaSSsyRdiHvj9cgRojKTB4esLYPs3YUsIpS6vK53bSvfJ
44SuvSX27wRsPNqUGridKT8l8MwEkfVgoQOfhmHnDL1MRUGeVmCs7Ug2P624+6n6
tM8J5yfs54IdQH+aDfzMYI58suPnYPymZPpwOIgtWsX8r9fg8nGjilmhzsAlNI0r
d8W1MsyUEZtqImw64LpWMyac94viyn6F9Vf3f3I7mzU6pE2lL3/F8eplIysBnGvM
EUmZjbJouqsGmmPBqXWqCt3kkooOS1mS1RnK3Dzdq0VNX2YYVjHHz4kW1j03igoG
a4Onw+tlyL0mLYq7XG36jvSbEHoqKJoY6MobZOZ2gKcVSeNA9WykuQ2rgQJImpbX
jMcuq4mlWOFObcm/s4kSPRw7mEmJ+NmxpmUus4LrI1E04Ts9U9gDcutT9BC9hC2T
VdEhVZLeEq3+dQ5mrAcz0mn6WrRca4/XJKCUPEKA+MNsdNxPDhfxO6mVi8uF+5br
dfiGmhUeW388qleXlDZeiLt7gh6uTOH+8ymCJlLQPWM/Qtv+iH4/Kzwge6Uiopim
DPq5cMTLqTdILSRzZNeidVJ0+UmfgCH2wakbFGHQ++TLxhhfgPePCaufqhC4njze
CkTd2lkZt+oMtBcG6u2Ejmu/gqPd4ejkQ58I16QK+ou/cqWLVCiijFb2RDNecdnj
csSmWwMdl0TnVUs8CfnoMLigHmkdnSASCnCbKeu0I0WwYPA6lbdPhgXVeU0qdBpj
BW+0Cp8FGEw7FCj/B+crk41qEe08z3CCV5olsuclvMF4+qidu+cpu9otNqYniz62
mCXegdb+h+NYbj4Rhcojx1/j3uKRgn0ldj6KJF3aKgDo6xeyIsM9j9ljGSAMGcVA
mzfqE0jT197qcVowuyu6G2KECSYqqAVmBzRhv2j41kSCVpEKa1hNd5JnD0UF1BqB
mYR0dKmnjbqwXBAqI4C8I9H2CBPqEUiLebXVBVb7sXkMcyY3/QwKpNWIFw98uvcr
ybWQ+du07QGm/FfXxKe+9JHiCxU24Z2DL+yA6zs9BnOpbEaEOPqZvvA7JH2EkJ3U
ZpbdqKgEtPfcBwklPaHWh9oUqmUTE/E35iZ1YQCW6LQsYlXuRS+yjiNV/vKqLQP8
s9SUrjTzh5EI3iUkJkZ4h00zJ0pFR3Xb7yLU0dhrXEVr/BN1MeRsIOQezK7fHrLG
FCq+cAi45cwHBvKfg73gqKete2LQoL9aJFHEoO6CZojDQLSLOV103U+UqxxSk8Wa
rja6lZcidUJN+E2Ce8QIPnGCqx1fn5S5phibZO40+HtE4b4lNAp9MWTQFrDfLT+i
XgONRfDTGlNYqT47bGY3pvHMVT0mxrRfT4g1HYSCPIUIFFo+1/F32zidgVHxM5/R
RHNfmQ1xM4cgOMRfhhl5PtHFAWsCeEBaqpwpSl4bug+bDnhXzAcLSsOwKSGAbyfr
pWGRV8x9EwuG/4j621A+xi6cl5/mnamlDg6qWTp8wUqw5GIF90dJ0MSs2TJjB3Vi
1iQUtef/GGw4wZIsq9Mug+VGfAYgqTeUN1o0rdV+GfxyY8h9g1b0gbqZddFRjMK7
2RmTQZLKRn48oryHDQf4Cezdef++U+nDNdqU/rnEwL0kG9RpANPjiefpkXQ8HMWx
XeopwERJT+F9n9r2YCSP7kXuTBpbEgfqmxJ2jh4Dx8eTfmKYINUwmeQoINyTY27W
+0bxsJq89Ipi4v8va4lKFbiSJtzFVSvylmDUYsPBCj1K/zyQKMcxJz9KU2jzeK/U
+ylTrUotWnb4ySt5jmdRZ8yIsrkOJ2aJYZNVnBUmzDEtY5FsSyFBYMrVYln0UgnU
XJMevVK8BnkAkY56Po5cVNsnAkpAJ6uoqsntzw3vLMobsPUeOhVLISnAJcEMcnDi
i9jCW3UEsYAwm8AdEh8WHBuZY4oD19d+NA8+LFcg+KNs70KbDnzIM+IGBqUorXUo
I2xa+/Px21aFFHKZYyLq9yvD+/wX7ig8Ke/7DOhwzsVzc0H1oCEzzlOvb0W3h+wK
0fI4gv3Rsfqg/XyvwGydoAoPunvVcf/dJ8TQHlomZVVgDfnfmYXcDb0+T6gciOUN
KLTaYXpoDJN+GuwZe3ZBcp5M4R7ZY7yaLe7LfZfcC+7nEpkxoesfJZPRpV0usNza
tYkz6ezifuftUq2411PCdT/G8nxZVwXdspeaT6bdYxpwl6HpFq9BL9O9HJ7kKBum
/zpy/iiubHSaWrztEPuUUyfUsNGhX1sHeOfm2UR/D370UZWviqyVq0BkomA9VjUM
aBg6m91k5ZvZ2P8VTYuzeTuri7rFa8KMUjz2SKtG+PdB9aLdPCce4C8VkBM4+2Dl
zdR3ht238mx50rCyXhm6zpF40bWvT3q1aKUp9vFBlPv061D1gsRh526KcQfdjvbo
T2VLnhm1XZb8sgBFJZRKWGDA1vE3B02ODNmGZX2mSxZxFJFDwhJZ/oa8jJ8KGsry
/Bk28se7LjzYAlytrZudR3TwL8aEHpxLQ416UR9hJdw3zZTelm7SRfAxbQKfIGoc
meaDr+WR0fn+hk/DbwWt0qHh9FP3FhQ0XrX1sdlMSyC7PLnCE8Z0OmhM01VYmbVM
PYE+z2pEd/eqZtFveRKfhbbCL4l8032vRiwY70LJPEmJbejiz3kssWLLfEqwN2Yc
tc9k69NYyj1uv9B/jZBCJExKDxbL/4oOSNQFsumSbEpnsnMiSda+1qp74qdYPRnR
OS9EEUjZRAvuysmt76sD+dvss18ibYxJ4Njfb0TTDVMo+MzPTCL0NVBtQWqXlwi3
cVVUfO1P9mDHo134AYB6dj137yODNnkvBMvAZ6oSNQusDXJfBve9UMdT94BYsf39
mRs+0CXvpsAT+GTQrevnTviOAOcj4YdWwiomzUEBBNLGEHL2JnXqoLUA8pz3yHLt
fFL7Y3cz7aXi2yR+6ciOaFMiZzZWIC3yacE3rfvS5Wgqi4eANZCylUcGLXj+VZkC
faClHWXYH/7wQKXdcColyZ9nG8iwfnWNRYh61kklIhsIreXxB+afwrl6zD1mn6y1
EIXSfbScC6/QGtzKwjFf0+f2vQlfP+L/I4oZ2eZ1qG+HoPZ+xMwyAVhCxLB2cjb9
xakOmt/b/zzysakNmZOEdeQLPougBO95fsh7YG/Awj4tOMOwqbNRMCRWJJVCeHwl
8MbK9IPh5WZ43OiCg4QVdDCDq/Qzpy6ql2D8wqKE8PRSWlH5PH4SWpnT9lBiB/tr
Bu/aogB205/929q4RM0RrdofaIQuZW/CPRfTD0yVK2UXGUPE5XmDM4m2wIQKrv1l
UogtDGUkiFdmYfXHNTmWodkGBZKYt514LeGRdNco9yr+cHkMbUCUCj0EhXHGGQDn
uoO06d2lEWFl3nRtCqNfle+5Mm/Rm+52TZhB/4E0+XdqHaN05SubKIclA3XKxGWA
uQoBFC63LfpVM+L4o6bIss8BR1WsPKponLCAV3ajZiDnzQUZ4c0zotS8CqWlxpSa
qxvNmisr9I12Nh+C5JmqLMz/Gl1PW7k3qUtyGhSPbxRWGDPSEx4Tk0RYMp1BDHXJ
8/0DqUzc4WynUdCiuSGfxj3Hiy4mJZbtHHKCjAxHa3GHrTaJIUENHTjXa9/T8fcT
6NhhT/Lz+gndpXOozFpRsrCKpsgphLsRWLn+bCato5W61Gjg8nC3ra1Ms7KzriFk
x/3wAAzl4Y1JVvdCkqkftOU7oim8ggJeF3ogH7glfkE2zZDsGb/RKrbkeOwStPyy
aMzJ6aV234/3S5fBUIAlw4ddJuP1ICFHN50GEdcY+aHJXHMqUfTrjnmqfXw9tuJH
wcljaZNWMLg+KRLI72+ucODPWZ6dGw/oHpELRodZNeyqgYOmlHjI3l/18CWCFEFA
EjDJEgOyNx+ILxQZmxb5NTIP1bNjPMAILSeoKfSDnXF9zvohLSjdZgUI+b7Jptu9
fUtmmzoteJ+uKz46u3JGqGO0NKdYS3T2okS9bLOO3qQsOxbSnd21wazhu81kYgzj
m0u8vMXbd2SrPin48NmnICGBbe/x0XXM9c1tMR6Q1A9SSlkPErKvUQbJfdL/c9/M
t1RAe94KT7CfJD0hztKYTNeTsS+z68Ti7rd111zR3xk/38xrjs4euV8GDQ7hmfje
aBPao1mZj0baqFNI5v3f52gS5QW/tH3NPFZuVFWllzzagdRKxgsa8iDja1JDvHsI
FNVWPy/UIYlEDZqxFxwQ4StJlAfi4bnrSzgTcSI355XNXfxJAV0gkzgQme89pXSX
t5/+/PLydPCe7nvebOfaOq+zeR77+Ebda/t2W9xxj5hLnkx26+TRNbz3kOfxg0Bd
36rHbuRqAAmxXNuH9vEKjp0G/5MapuadfRdiwZCKXOTOELy0qlCTc6AiBRYbOAqI
pVDm7w6SrlcrF5tRYeqC0gUsAYf1ANCBCot82MlJqYrdAtS1sULLS/KrB1Mlml0J
ITzsjpQ0O2jbf9+gXstPnEObKJhwEk6uPsCOwHxXhofxQG/lCSS1TGrNgpNPJ8+o
GLDfXrrdy2WUXcV9HM2S6ODPujg0eGlRe7wg1N4PeJtD7N0BCMnHMB6AUNDNcQir
smtaIvAZMLjCehSLLTf2EPbFg9+zp5hKZEooRmKCvPG9aGr/GhHbzZDQ2t8qraB3
Ma6angmYK5OO/sM6+Ok5PjmXVOS+2hDh3XTFwJqsksGhX0AkrtKeB3dLZwVGQWoj
7YRNmhqbXMA8jXjTMdAWka1bq+nPoDjE6FTqq4/WjvZKUGGn8+sDI21IAfywm5Nr
pu4vNNodxtMhWrl88o+EcVsoYb5Zk3HROeovxfNgDNgASH8pwjPdI4aV6YH5bakj
0L6+AzO0vYc136mQjGjqTGyWhM7/f0iMf+Tz9MUasTDjS3znpOVvtVt40tA+ZTOz
QJRKhiXWiM1jeYYVG6gFlRURN81IE1g4J4ITdweahC1t2nib9Hz0X/fdD2LTme26
L6357bocAmZ3otf+YvwTQOVHNTl7EXXlDCdA1IGHhp1Y/949DXIC7Y38ldyH5GZV
Rzu2/vTZ74eTS0JctmtQr1gyEOdo1F/dQD06+E19bF61bZ0/BBFcyi3Q3i/4M6nv
BaBO1Xr2DqJYW6y5JuNUDukCKr6cxLaZyI2WBSQfsmpr+kPo9TZK/wyJB1TNJYf0
ukTcUp5LYILCBjPPm/8RXSnN6d7D8nCWvtCPsZJMBZ6DqVH4p9rrKskYeBC0qzIu
UW9QzH+esQAo/qqndZ6d0s53rIgAkWrfv9P5QSJkPzrw4cZEXU95+YD3Yqs0kLk4
7ftn1rqw9CfjKt6cE35KVBMH8C6z/6MBWHFo+qyUMQFfzhXym+ySbT4YqdHFoxwu
uhdCHKmVmlCjSGHgcaQ/8B9bpiGqYXtEhIqIonILP2yYyoYuiQihYsepcJegJ8zd
XKaOiKC9yqYUIoDNnMlZNhWiYRK2dpIBm5bxyC98G3IZN+fbuihvh5Q7yPCv80Gq
iSIYU92OkqTt/o/EU9rgRbl+dmh8vYv2A4yqUXJP2xg2Rg51v1jt2wLG5CPl6hyD
0isdaL7nj4vCIlt5HCqIvqLd/sl7eL15Y4B8bUXdPbdKBczjhoVG8V3IYAvpy6lX
vyhQ4dSWh8cdfmy0RMp0WyRGucOGoZgNHDFUYThHhWEI7cmAahnOZcti4ngKNUp8
Sxr/Lm3aQKchfTacTD3tssIFr1M1Z7xgwFmUW5YZKSQfJUIknJR0qZoXdgcacEeu
WhoRSO/9i67QwqtfwLQ6vj6ziQ19tEYKwDpQBRYWFPBDF2NThINFLcwp8DsvTaJj
P2tdUtyey+hJ3FkGPdfbRnqBBwWYHkB0Bmw6utD0fx+ZVR4RxXuQNAXAR7UApkED
LXYNCq9z/Fw9IrQ6xOCK9bYwETKjsba/L9T5oScyaPaaNM5vGCTjCa0knoVOW2d0
WGA8aBHWrWqUkO5+v10IvMbn/8UqGryYftnCdxsSqGUL93eAVJmKTwYDMm/UNu5Y
vwWyXsjTwyj533w6aVHpJCy+C2QWTzyBk1TpDAWYjzfXo/v33tu4Ng3ZYgqOh7sl
1etvSReBYdhzMXzMXKQ3q2MKMmsQwcgRxXvo6AZtjBBfa164eYImy9FePjjkVvQp
ifZd03dyncPSgivk4gKKSXqB5+cyKiODGZW2Th8ENwquUUaAZnQXUi460qIP84u8
pBn9rbsCxjlf4/FzS2H1JwechhfEpTgmICu8WPyCGNd0NuwOBAkvmZgkcRD7uBMq
hKjWz22Cw4s931rRtRcWMohJtsDfeagI9h4RiH+8zZxOQDg/2FqU8hElhMP1P6Vi
MzIfYCGbX720LJ8GDdAehRdb+r3tPxkltaPQbFwgXfSrmFf86Dx5rfjFR7jJSThF
`pragma protect end_protected
